
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"e7",x"fe",x"49",x"72"),
     1 => (x"9a",x"4a",x"13",x"87"),
     2 => (x"fe",x"87",x"f5",x"05"),
     3 => (x"c2",x"1e",x"87",x"da"),
     4 => (x"49",x"bf",x"cd",x"f6"),
     5 => (x"48",x"cd",x"f6",x"c2"),
     6 => (x"c4",x"78",x"a1",x"c1"),
     7 => (x"03",x"a9",x"b7",x"c0"),
     8 => (x"d4",x"ff",x"87",x"db"),
     9 => (x"d1",x"f6",x"c2",x"48"),
    10 => (x"f6",x"c2",x"78",x"bf"),
    11 => (x"c2",x"49",x"bf",x"cd"),
    12 => (x"c1",x"48",x"cd",x"f6"),
    13 => (x"c0",x"c4",x"78",x"a1"),
    14 => (x"e5",x"04",x"a9",x"b7"),
    15 => (x"48",x"d0",x"ff",x"87"),
    16 => (x"f6",x"c2",x"78",x"c8"),
    17 => (x"78",x"c0",x"48",x"d9"),
    18 => (x"00",x"00",x"4f",x"26"),
    19 => (x"00",x"00",x"00",x"00"),
    20 => (x"00",x"00",x"00",x"00"),
    21 => (x"00",x"5f",x"5f",x"00"),
    22 => (x"03",x"00",x"00",x"00"),
    23 => (x"03",x"03",x"00",x"03"),
    24 => (x"7f",x"14",x"00",x"00"),
    25 => (x"7f",x"7f",x"14",x"7f"),
    26 => (x"24",x"00",x"00",x"14"),
    27 => (x"3a",x"6b",x"6b",x"2e"),
    28 => (x"6a",x"4c",x"00",x"12"),
    29 => (x"56",x"6c",x"18",x"36"),
    30 => (x"7e",x"30",x"00",x"32"),
    31 => (x"3a",x"77",x"59",x"4f"),
    32 => (x"00",x"00",x"40",x"68"),
    33 => (x"00",x"03",x"07",x"04"),
    34 => (x"00",x"00",x"00",x"00"),
    35 => (x"41",x"63",x"3e",x"1c"),
    36 => (x"00",x"00",x"00",x"00"),
    37 => (x"1c",x"3e",x"63",x"41"),
    38 => (x"2a",x"08",x"00",x"00"),
    39 => (x"3e",x"1c",x"1c",x"3e"),
    40 => (x"08",x"00",x"08",x"2a"),
    41 => (x"08",x"3e",x"3e",x"08"),
    42 => (x"00",x"00",x"00",x"08"),
    43 => (x"00",x"60",x"e0",x"80"),
    44 => (x"08",x"00",x"00",x"00"),
    45 => (x"08",x"08",x"08",x"08"),
    46 => (x"00",x"00",x"00",x"08"),
    47 => (x"00",x"60",x"60",x"00"),
    48 => (x"60",x"40",x"00",x"00"),
    49 => (x"06",x"0c",x"18",x"30"),
    50 => (x"3e",x"00",x"01",x"03"),
    51 => (x"7f",x"4d",x"59",x"7f"),
    52 => (x"04",x"00",x"00",x"3e"),
    53 => (x"00",x"7f",x"7f",x"06"),
    54 => (x"42",x"00",x"00",x"00"),
    55 => (x"4f",x"59",x"71",x"63"),
    56 => (x"22",x"00",x"00",x"46"),
    57 => (x"7f",x"49",x"49",x"63"),
    58 => (x"1c",x"18",x"00",x"36"),
    59 => (x"7f",x"7f",x"13",x"16"),
    60 => (x"27",x"00",x"00",x"10"),
    61 => (x"7d",x"45",x"45",x"67"),
    62 => (x"3c",x"00",x"00",x"39"),
    63 => (x"79",x"49",x"4b",x"7e"),
    64 => (x"01",x"00",x"00",x"30"),
    65 => (x"0f",x"79",x"71",x"01"),
    66 => (x"36",x"00",x"00",x"07"),
    67 => (x"7f",x"49",x"49",x"7f"),
    68 => (x"06",x"00",x"00",x"36"),
    69 => (x"3f",x"69",x"49",x"4f"),
    70 => (x"00",x"00",x"00",x"1e"),
    71 => (x"00",x"66",x"66",x"00"),
    72 => (x"00",x"00",x"00",x"00"),
    73 => (x"00",x"66",x"e6",x"80"),
    74 => (x"08",x"00",x"00",x"00"),
    75 => (x"22",x"14",x"14",x"08"),
    76 => (x"14",x"00",x"00",x"22"),
    77 => (x"14",x"14",x"14",x"14"),
    78 => (x"22",x"00",x"00",x"14"),
    79 => (x"08",x"14",x"14",x"22"),
    80 => (x"02",x"00",x"00",x"08"),
    81 => (x"0f",x"59",x"51",x"03"),
    82 => (x"7f",x"3e",x"00",x"06"),
    83 => (x"1f",x"55",x"5d",x"41"),
    84 => (x"7e",x"00",x"00",x"1e"),
    85 => (x"7f",x"09",x"09",x"7f"),
    86 => (x"7f",x"00",x"00",x"7e"),
    87 => (x"7f",x"49",x"49",x"7f"),
    88 => (x"1c",x"00",x"00",x"36"),
    89 => (x"41",x"41",x"63",x"3e"),
    90 => (x"7f",x"00",x"00",x"41"),
    91 => (x"3e",x"63",x"41",x"7f"),
    92 => (x"7f",x"00",x"00",x"1c"),
    93 => (x"41",x"49",x"49",x"7f"),
    94 => (x"7f",x"00",x"00",x"41"),
    95 => (x"01",x"09",x"09",x"7f"),
    96 => (x"3e",x"00",x"00",x"01"),
    97 => (x"7b",x"49",x"41",x"7f"),
    98 => (x"7f",x"00",x"00",x"7a"),
    99 => (x"7f",x"08",x"08",x"7f"),
   100 => (x"00",x"00",x"00",x"7f"),
   101 => (x"41",x"7f",x"7f",x"41"),
   102 => (x"20",x"00",x"00",x"00"),
   103 => (x"7f",x"40",x"40",x"60"),
   104 => (x"7f",x"7f",x"00",x"3f"),
   105 => (x"63",x"36",x"1c",x"08"),
   106 => (x"7f",x"00",x"00",x"41"),
   107 => (x"40",x"40",x"40",x"7f"),
   108 => (x"7f",x"7f",x"00",x"40"),
   109 => (x"7f",x"06",x"0c",x"06"),
   110 => (x"7f",x"7f",x"00",x"7f"),
   111 => (x"7f",x"18",x"0c",x"06"),
   112 => (x"3e",x"00",x"00",x"7f"),
   113 => (x"7f",x"41",x"41",x"7f"),
   114 => (x"7f",x"00",x"00",x"3e"),
   115 => (x"0f",x"09",x"09",x"7f"),
   116 => (x"7f",x"3e",x"00",x"06"),
   117 => (x"7e",x"7f",x"61",x"41"),
   118 => (x"7f",x"00",x"00",x"40"),
   119 => (x"7f",x"19",x"09",x"7f"),
   120 => (x"26",x"00",x"00",x"66"),
   121 => (x"7b",x"59",x"4d",x"6f"),
   122 => (x"01",x"00",x"00",x"32"),
   123 => (x"01",x"7f",x"7f",x"01"),
   124 => (x"3f",x"00",x"00",x"01"),
   125 => (x"7f",x"40",x"40",x"7f"),
   126 => (x"0f",x"00",x"00",x"3f"),
   127 => (x"3f",x"70",x"70",x"3f"),
   128 => (x"7f",x"7f",x"00",x"0f"),
   129 => (x"7f",x"30",x"18",x"30"),
   130 => (x"63",x"41",x"00",x"7f"),
   131 => (x"36",x"1c",x"1c",x"36"),
   132 => (x"03",x"01",x"41",x"63"),
   133 => (x"06",x"7c",x"7c",x"06"),
   134 => (x"71",x"61",x"01",x"03"),
   135 => (x"43",x"47",x"4d",x"59"),
   136 => (x"00",x"00",x"00",x"41"),
   137 => (x"41",x"41",x"7f",x"7f"),
   138 => (x"03",x"01",x"00",x"00"),
   139 => (x"30",x"18",x"0c",x"06"),
   140 => (x"00",x"00",x"40",x"60"),
   141 => (x"7f",x"7f",x"41",x"41"),
   142 => (x"0c",x"08",x"00",x"00"),
   143 => (x"0c",x"06",x"03",x"06"),
   144 => (x"80",x"80",x"00",x"08"),
   145 => (x"80",x"80",x"80",x"80"),
   146 => (x"00",x"00",x"00",x"80"),
   147 => (x"04",x"07",x"03",x"00"),
   148 => (x"20",x"00",x"00",x"00"),
   149 => (x"7c",x"54",x"54",x"74"),
   150 => (x"7f",x"00",x"00",x"78"),
   151 => (x"7c",x"44",x"44",x"7f"),
   152 => (x"38",x"00",x"00",x"38"),
   153 => (x"44",x"44",x"44",x"7c"),
   154 => (x"38",x"00",x"00",x"00"),
   155 => (x"7f",x"44",x"44",x"7c"),
   156 => (x"38",x"00",x"00",x"7f"),
   157 => (x"5c",x"54",x"54",x"7c"),
   158 => (x"04",x"00",x"00",x"18"),
   159 => (x"05",x"05",x"7f",x"7e"),
   160 => (x"18",x"00",x"00",x"00"),
   161 => (x"fc",x"a4",x"a4",x"bc"),
   162 => (x"7f",x"00",x"00",x"7c"),
   163 => (x"7c",x"04",x"04",x"7f"),
   164 => (x"00",x"00",x"00",x"78"),
   165 => (x"40",x"7d",x"3d",x"00"),
   166 => (x"80",x"00",x"00",x"00"),
   167 => (x"7d",x"fd",x"80",x"80"),
   168 => (x"7f",x"00",x"00",x"00"),
   169 => (x"6c",x"38",x"10",x"7f"),
   170 => (x"00",x"00",x"00",x"44"),
   171 => (x"40",x"7f",x"3f",x"00"),
   172 => (x"7c",x"7c",x"00",x"00"),
   173 => (x"7c",x"0c",x"18",x"0c"),
   174 => (x"7c",x"00",x"00",x"78"),
   175 => (x"7c",x"04",x"04",x"7c"),
   176 => (x"38",x"00",x"00",x"78"),
   177 => (x"7c",x"44",x"44",x"7c"),
   178 => (x"fc",x"00",x"00",x"38"),
   179 => (x"3c",x"24",x"24",x"fc"),
   180 => (x"18",x"00",x"00",x"18"),
   181 => (x"fc",x"24",x"24",x"3c"),
   182 => (x"7c",x"00",x"00",x"fc"),
   183 => (x"0c",x"04",x"04",x"7c"),
   184 => (x"48",x"00",x"00",x"08"),
   185 => (x"74",x"54",x"54",x"5c"),
   186 => (x"04",x"00",x"00",x"20"),
   187 => (x"44",x"44",x"7f",x"3f"),
   188 => (x"3c",x"00",x"00",x"00"),
   189 => (x"7c",x"40",x"40",x"7c"),
   190 => (x"1c",x"00",x"00",x"7c"),
   191 => (x"3c",x"60",x"60",x"3c"),
   192 => (x"7c",x"3c",x"00",x"1c"),
   193 => (x"7c",x"60",x"30",x"60"),
   194 => (x"6c",x"44",x"00",x"3c"),
   195 => (x"6c",x"38",x"10",x"38"),
   196 => (x"1c",x"00",x"00",x"44"),
   197 => (x"3c",x"60",x"e0",x"bc"),
   198 => (x"44",x"00",x"00",x"1c"),
   199 => (x"4c",x"5c",x"74",x"64"),
   200 => (x"08",x"00",x"00",x"44"),
   201 => (x"41",x"77",x"3e",x"08"),
   202 => (x"00",x"00",x"00",x"41"),
   203 => (x"00",x"7f",x"7f",x"00"),
   204 => (x"41",x"00",x"00",x"00"),
   205 => (x"08",x"3e",x"77",x"41"),
   206 => (x"01",x"02",x"00",x"08"),
   207 => (x"02",x"02",x"03",x"01"),
   208 => (x"7f",x"7f",x"00",x"01"),
   209 => (x"7f",x"7f",x"7f",x"7f"),
   210 => (x"08",x"08",x"00",x"7f"),
   211 => (x"3e",x"3e",x"1c",x"1c"),
   212 => (x"7f",x"7f",x"7f",x"7f"),
   213 => (x"1c",x"1c",x"3e",x"3e"),
   214 => (x"10",x"00",x"08",x"08"),
   215 => (x"18",x"7c",x"7c",x"18"),
   216 => (x"10",x"00",x"00",x"10"),
   217 => (x"30",x"7c",x"7c",x"30"),
   218 => (x"30",x"10",x"00",x"10"),
   219 => (x"1e",x"78",x"60",x"60"),
   220 => (x"66",x"42",x"00",x"06"),
   221 => (x"66",x"3c",x"18",x"3c"),
   222 => (x"38",x"78",x"00",x"42"),
   223 => (x"6c",x"c6",x"c2",x"6a"),
   224 => (x"00",x"60",x"00",x"38"),
   225 => (x"00",x"00",x"60",x"00"),
   226 => (x"5e",x"0e",x"00",x"60"),
   227 => (x"0e",x"5d",x"5c",x"5b"),
   228 => (x"c2",x"4c",x"71",x"1e"),
   229 => (x"4d",x"bf",x"ea",x"f6"),
   230 => (x"1e",x"c0",x"4b",x"c0"),
   231 => (x"c7",x"02",x"ab",x"74"),
   232 => (x"48",x"a6",x"c4",x"87"),
   233 => (x"87",x"c5",x"78",x"c0"),
   234 => (x"c1",x"48",x"a6",x"c4"),
   235 => (x"1e",x"66",x"c4",x"78"),
   236 => (x"df",x"ee",x"49",x"73"),
   237 => (x"c0",x"86",x"c8",x"87"),
   238 => (x"ef",x"ef",x"49",x"e0"),
   239 => (x"4a",x"a5",x"c4",x"87"),
   240 => (x"f0",x"f0",x"49",x"6a"),
   241 => (x"87",x"c6",x"f1",x"87"),
   242 => (x"83",x"c1",x"85",x"cb"),
   243 => (x"04",x"ab",x"b7",x"c8"),
   244 => (x"26",x"87",x"c7",x"ff"),
   245 => (x"4c",x"26",x"4d",x"26"),
   246 => (x"4f",x"26",x"4b",x"26"),
   247 => (x"c2",x"4a",x"71",x"1e"),
   248 => (x"c2",x"5a",x"ee",x"f6"),
   249 => (x"c7",x"48",x"ee",x"f6"),
   250 => (x"dd",x"fe",x"49",x"78"),
   251 => (x"1e",x"4f",x"26",x"87"),
   252 => (x"4a",x"71",x"1e",x"73"),
   253 => (x"03",x"aa",x"b7",x"c0"),
   254 => (x"dd",x"c2",x"87",x"d3"),
   255 => (x"c4",x"05",x"bf",x"cf"),
   256 => (x"c2",x"4b",x"c1",x"87"),
   257 => (x"c2",x"4b",x"c0",x"87"),
   258 => (x"c4",x"5b",x"d3",x"dd"),
   259 => (x"d3",x"dd",x"c2",x"87"),
   260 => (x"cf",x"dd",x"c2",x"5a"),
   261 => (x"9a",x"c1",x"4a",x"bf"),
   262 => (x"49",x"a2",x"c0",x"c1"),
   263 => (x"fc",x"87",x"e8",x"ec"),
   264 => (x"cf",x"dd",x"c2",x"48"),
   265 => (x"ef",x"fe",x"78",x"bf"),
   266 => (x"4a",x"71",x"1e",x"87"),
   267 => (x"72",x"1e",x"66",x"c4"),
   268 => (x"da",x"df",x"ff",x"49"),
   269 => (x"4f",x"26",x"26",x"87"),
   270 => (x"cf",x"dd",x"c2",x"1e"),
   271 => (x"dc",x"ff",x"49",x"bf"),
   272 => (x"f6",x"c2",x"87",x"c2"),
   273 => (x"bf",x"e8",x"48",x"e2"),
   274 => (x"de",x"f6",x"c2",x"78"),
   275 => (x"78",x"bf",x"ec",x"48"),
   276 => (x"bf",x"e2",x"f6",x"c2"),
   277 => (x"ff",x"c3",x"49",x"4a"),
   278 => (x"2a",x"b7",x"c8",x"99"),
   279 => (x"b0",x"71",x"48",x"72"),
   280 => (x"58",x"ea",x"f6",x"c2"),
   281 => (x"5e",x"0e",x"4f",x"26"),
   282 => (x"0e",x"5d",x"5c",x"5b"),
   283 => (x"c7",x"ff",x"4b",x"71"),
   284 => (x"dd",x"f6",x"c2",x"87"),
   285 => (x"73",x"50",x"c0",x"48"),
   286 => (x"e7",x"db",x"ff",x"49"),
   287 => (x"4c",x"49",x"70",x"87"),
   288 => (x"ee",x"cb",x"9c",x"c2"),
   289 => (x"87",x"cf",x"cb",x"49"),
   290 => (x"c2",x"4d",x"49",x"70"),
   291 => (x"bf",x"97",x"dd",x"f6"),
   292 => (x"87",x"e4",x"c1",x"05"),
   293 => (x"c2",x"49",x"66",x"d0"),
   294 => (x"99",x"bf",x"e6",x"f6"),
   295 => (x"d4",x"87",x"d7",x"05"),
   296 => (x"f6",x"c2",x"49",x"66"),
   297 => (x"05",x"99",x"bf",x"de"),
   298 => (x"49",x"73",x"87",x"cc"),
   299 => (x"87",x"f4",x"da",x"ff"),
   300 => (x"c1",x"02",x"98",x"70"),
   301 => (x"4c",x"c1",x"87",x"c2"),
   302 => (x"75",x"87",x"fd",x"fd"),
   303 => (x"87",x"e3",x"ca",x"49"),
   304 => (x"c6",x"02",x"98",x"70"),
   305 => (x"dd",x"f6",x"c2",x"87"),
   306 => (x"c2",x"50",x"c1",x"48"),
   307 => (x"bf",x"97",x"dd",x"f6"),
   308 => (x"87",x"e4",x"c0",x"05"),
   309 => (x"bf",x"e6",x"f6",x"c2"),
   310 => (x"99",x"66",x"d0",x"49"),
   311 => (x"87",x"d6",x"ff",x"05"),
   312 => (x"bf",x"de",x"f6",x"c2"),
   313 => (x"99",x"66",x"d4",x"49"),
   314 => (x"87",x"ca",x"ff",x"05"),
   315 => (x"d9",x"ff",x"49",x"73"),
   316 => (x"98",x"70",x"87",x"f2"),
   317 => (x"87",x"fe",x"fe",x"05"),
   318 => (x"d7",x"fb",x"48",x"74"),
   319 => (x"5b",x"5e",x"0e",x"87"),
   320 => (x"f4",x"0e",x"5d",x"5c"),
   321 => (x"4c",x"4d",x"c0",x"86"),
   322 => (x"c4",x"7e",x"bf",x"ec"),
   323 => (x"f6",x"c2",x"48",x"a6"),
   324 => (x"c1",x"78",x"bf",x"ea"),
   325 => (x"c7",x"1e",x"c0",x"1e"),
   326 => (x"87",x"ca",x"fd",x"49"),
   327 => (x"98",x"70",x"86",x"c8"),
   328 => (x"ff",x"87",x"ce",x"02"),
   329 => (x"87",x"c7",x"fb",x"49"),
   330 => (x"ff",x"49",x"da",x"c1"),
   331 => (x"c1",x"87",x"f5",x"d8"),
   332 => (x"dd",x"f6",x"c2",x"4d"),
   333 => (x"c3",x"02",x"bf",x"97"),
   334 => (x"87",x"f9",x"cd",x"87"),
   335 => (x"bf",x"e2",x"f6",x"c2"),
   336 => (x"cf",x"dd",x"c2",x"4b"),
   337 => (x"eb",x"c0",x"05",x"bf"),
   338 => (x"49",x"fd",x"c3",x"87"),
   339 => (x"87",x"d4",x"d8",x"ff"),
   340 => (x"ff",x"49",x"fa",x"c3"),
   341 => (x"73",x"87",x"cd",x"d8"),
   342 => (x"99",x"ff",x"c3",x"49"),
   343 => (x"49",x"c0",x"1e",x"71"),
   344 => (x"73",x"87",x"c6",x"fb"),
   345 => (x"29",x"b7",x"c8",x"49"),
   346 => (x"49",x"c1",x"1e",x"71"),
   347 => (x"c8",x"87",x"fa",x"fa"),
   348 => (x"87",x"c1",x"c6",x"86"),
   349 => (x"bf",x"e6",x"f6",x"c2"),
   350 => (x"dd",x"02",x"9b",x"4b"),
   351 => (x"cb",x"dd",x"c2",x"87"),
   352 => (x"de",x"c7",x"49",x"bf"),
   353 => (x"05",x"98",x"70",x"87"),
   354 => (x"4b",x"c0",x"87",x"c4"),
   355 => (x"e0",x"c2",x"87",x"d2"),
   356 => (x"87",x"c3",x"c7",x"49"),
   357 => (x"58",x"cf",x"dd",x"c2"),
   358 => (x"dd",x"c2",x"87",x"c6"),
   359 => (x"78",x"c0",x"48",x"cb"),
   360 => (x"99",x"c2",x"49",x"73"),
   361 => (x"c3",x"87",x"ce",x"05"),
   362 => (x"d6",x"ff",x"49",x"eb"),
   363 => (x"49",x"70",x"87",x"f6"),
   364 => (x"c2",x"02",x"99",x"c2"),
   365 => (x"73",x"4c",x"fb",x"87"),
   366 => (x"05",x"99",x"c1",x"49"),
   367 => (x"f4",x"c3",x"87",x"ce"),
   368 => (x"df",x"d6",x"ff",x"49"),
   369 => (x"c2",x"49",x"70",x"87"),
   370 => (x"87",x"c2",x"02",x"99"),
   371 => (x"49",x"73",x"4c",x"fa"),
   372 => (x"ce",x"05",x"99",x"c8"),
   373 => (x"49",x"f5",x"c3",x"87"),
   374 => (x"87",x"c8",x"d6",x"ff"),
   375 => (x"99",x"c2",x"49",x"70"),
   376 => (x"c2",x"87",x"d5",x"02"),
   377 => (x"02",x"bf",x"ee",x"f6"),
   378 => (x"c1",x"48",x"87",x"ca"),
   379 => (x"f2",x"f6",x"c2",x"88"),
   380 => (x"87",x"c2",x"c0",x"58"),
   381 => (x"4d",x"c1",x"4c",x"ff"),
   382 => (x"99",x"c4",x"49",x"73"),
   383 => (x"c3",x"87",x"ce",x"05"),
   384 => (x"d5",x"ff",x"49",x"f2"),
   385 => (x"49",x"70",x"87",x"de"),
   386 => (x"dc",x"02",x"99",x"c2"),
   387 => (x"ee",x"f6",x"c2",x"87"),
   388 => (x"c7",x"48",x"7e",x"bf"),
   389 => (x"c0",x"03",x"a8",x"b7"),
   390 => (x"48",x"6e",x"87",x"cb"),
   391 => (x"f6",x"c2",x"80",x"c1"),
   392 => (x"c2",x"c0",x"58",x"f2"),
   393 => (x"c1",x"4c",x"fe",x"87"),
   394 => (x"49",x"fd",x"c3",x"4d"),
   395 => (x"87",x"f4",x"d4",x"ff"),
   396 => (x"99",x"c2",x"49",x"70"),
   397 => (x"87",x"d5",x"c0",x"02"),
   398 => (x"bf",x"ee",x"f6",x"c2"),
   399 => (x"87",x"c9",x"c0",x"02"),
   400 => (x"48",x"ee",x"f6",x"c2"),
   401 => (x"c2",x"c0",x"78",x"c0"),
   402 => (x"c1",x"4c",x"fd",x"87"),
   403 => (x"49",x"fa",x"c3",x"4d"),
   404 => (x"87",x"d0",x"d4",x"ff"),
   405 => (x"99",x"c2",x"49",x"70"),
   406 => (x"87",x"d9",x"c0",x"02"),
   407 => (x"bf",x"ee",x"f6",x"c2"),
   408 => (x"a8",x"b7",x"c7",x"48"),
   409 => (x"87",x"c9",x"c0",x"03"),
   410 => (x"48",x"ee",x"f6",x"c2"),
   411 => (x"c2",x"c0",x"78",x"c7"),
   412 => (x"c1",x"4c",x"fc",x"87"),
   413 => (x"ac",x"b7",x"c0",x"4d"),
   414 => (x"87",x"d1",x"c0",x"03"),
   415 => (x"c1",x"4a",x"66",x"c4"),
   416 => (x"02",x"6a",x"82",x"d8"),
   417 => (x"6a",x"87",x"c6",x"c0"),
   418 => (x"73",x"49",x"74",x"4b"),
   419 => (x"c3",x"1e",x"c0",x"0f"),
   420 => (x"da",x"c1",x"1e",x"f0"),
   421 => (x"87",x"ce",x"f7",x"49"),
   422 => (x"98",x"70",x"86",x"c8"),
   423 => (x"87",x"e2",x"c0",x"02"),
   424 => (x"c2",x"48",x"a6",x"c8"),
   425 => (x"78",x"bf",x"ee",x"f6"),
   426 => (x"cb",x"49",x"66",x"c8"),
   427 => (x"48",x"66",x"c4",x"91"),
   428 => (x"7e",x"70",x"80",x"71"),
   429 => (x"c0",x"02",x"bf",x"6e"),
   430 => (x"bf",x"6e",x"87",x"c8"),
   431 => (x"49",x"66",x"c8",x"4b"),
   432 => (x"9d",x"75",x"0f",x"73"),
   433 => (x"87",x"c8",x"c0",x"02"),
   434 => (x"bf",x"ee",x"f6",x"c2"),
   435 => (x"87",x"fa",x"f2",x"49"),
   436 => (x"bf",x"d3",x"dd",x"c2"),
   437 => (x"87",x"dd",x"c0",x"02"),
   438 => (x"87",x"c7",x"c2",x"49"),
   439 => (x"c0",x"02",x"98",x"70"),
   440 => (x"f6",x"c2",x"87",x"d3"),
   441 => (x"f2",x"49",x"bf",x"ee"),
   442 => (x"49",x"c0",x"87",x"e0"),
   443 => (x"c2",x"87",x"c0",x"f4"),
   444 => (x"c0",x"48",x"d3",x"dd"),
   445 => (x"f3",x"8e",x"f4",x"78"),
   446 => (x"5e",x"0e",x"87",x"da"),
   447 => (x"0e",x"5d",x"5c",x"5b"),
   448 => (x"c2",x"4c",x"71",x"1e"),
   449 => (x"49",x"bf",x"ea",x"f6"),
   450 => (x"4d",x"a1",x"cd",x"c1"),
   451 => (x"69",x"81",x"d1",x"c1"),
   452 => (x"02",x"9c",x"74",x"7e"),
   453 => (x"a5",x"c4",x"87",x"cf"),
   454 => (x"c2",x"7b",x"74",x"4b"),
   455 => (x"49",x"bf",x"ea",x"f6"),
   456 => (x"6e",x"87",x"f9",x"f2"),
   457 => (x"05",x"9c",x"74",x"7b"),
   458 => (x"4b",x"c0",x"87",x"c4"),
   459 => (x"4b",x"c1",x"87",x"c2"),
   460 => (x"fa",x"f2",x"49",x"73"),
   461 => (x"02",x"66",x"d4",x"87"),
   462 => (x"da",x"49",x"87",x"c7"),
   463 => (x"c2",x"4a",x"70",x"87"),
   464 => (x"c2",x"4a",x"c0",x"87"),
   465 => (x"26",x"5a",x"d7",x"dd"),
   466 => (x"00",x"87",x"c9",x"f2"),
   467 => (x"00",x"00",x"00",x"00"),
   468 => (x"00",x"00",x"00",x"00"),
   469 => (x"1e",x"00",x"00",x"00"),
   470 => (x"c8",x"ff",x"4a",x"71"),
   471 => (x"a1",x"72",x"49",x"bf"),
   472 => (x"1e",x"4f",x"26",x"48"),
   473 => (x"89",x"bf",x"c8",x"ff"),
   474 => (x"c0",x"c0",x"c0",x"fe"),
   475 => (x"01",x"a9",x"c0",x"c0"),
   476 => (x"4a",x"c0",x"87",x"c4"),
   477 => (x"4a",x"c1",x"87",x"c2"),
   478 => (x"4f",x"26",x"48",x"72"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"71",x"1e",x"0e",x"5d"),
   481 => (x"4b",x"d4",x"ff",x"4d"),
   482 => (x"f6",x"c2",x"1e",x"75"),
   483 => (x"c1",x"fe",x"49",x"f2"),
   484 => (x"86",x"c4",x"87",x"d0"),
   485 => (x"02",x"6e",x"7e",x"70"),
   486 => (x"c2",x"87",x"ff",x"c3"),
   487 => (x"4c",x"bf",x"fa",x"f6"),
   488 => (x"da",x"fe",x"49",x"75"),
   489 => (x"a8",x"de",x"87",x"fe"),
   490 => (x"87",x"eb",x"c0",x"05"),
   491 => (x"d3",x"ff",x"49",x"75"),
   492 => (x"98",x"70",x"87",x"ec"),
   493 => (x"c2",x"87",x"db",x"02"),
   494 => (x"1e",x"bf",x"f5",x"f5"),
   495 => (x"ff",x"49",x"e1",x"c0"),
   496 => (x"c4",x"87",x"f7",x"d0"),
   497 => (x"f4",x"e2",x"c2",x"86"),
   498 => (x"c2",x"50",x"c0",x"48"),
   499 => (x"fe",x"49",x"c1",x"f6"),
   500 => (x"48",x"c1",x"87",x"ea"),
   501 => (x"ff",x"87",x"c5",x"c3"),
   502 => (x"c5",x"c8",x"48",x"d0"),
   503 => (x"7b",x"d6",x"c1",x"78"),
   504 => (x"97",x"6e",x"4a",x"c0"),
   505 => (x"48",x"6e",x"7b",x"bf"),
   506 => (x"7e",x"70",x"80",x"c1"),
   507 => (x"e0",x"c0",x"82",x"c1"),
   508 => (x"ff",x"04",x"aa",x"b7"),
   509 => (x"d0",x"ff",x"87",x"ec"),
   510 => (x"c8",x"78",x"c4",x"48"),
   511 => (x"d3",x"c1",x"78",x"c5"),
   512 => (x"c4",x"7b",x"c1",x"7b"),
   513 => (x"02",x"9c",x"74",x"78"),
   514 => (x"c2",x"87",x"fd",x"c1"),
   515 => (x"c8",x"7e",x"ee",x"e4"),
   516 => (x"c0",x"8c",x"4d",x"c0"),
   517 => (x"c6",x"03",x"ac",x"b7"),
   518 => (x"a4",x"c0",x"c8",x"87"),
   519 => (x"c2",x"4c",x"c0",x"4d"),
   520 => (x"bf",x"97",x"df",x"f1"),
   521 => (x"02",x"99",x"d0",x"49"),
   522 => (x"1e",x"c0",x"87",x"d2"),
   523 => (x"49",x"f2",x"f6",x"c2"),
   524 => (x"87",x"ca",x"c2",x"fe"),
   525 => (x"49",x"70",x"86",x"c4"),
   526 => (x"87",x"ef",x"c0",x"4a"),
   527 => (x"1e",x"ee",x"e4",x"c2"),
   528 => (x"49",x"f2",x"f6",x"c2"),
   529 => (x"87",x"f6",x"c1",x"fe"),
   530 => (x"49",x"70",x"86",x"c4"),
   531 => (x"48",x"d0",x"ff",x"4a"),
   532 => (x"c1",x"78",x"c5",x"c8"),
   533 => (x"97",x"6e",x"7b",x"d4"),
   534 => (x"48",x"6e",x"7b",x"bf"),
   535 => (x"7e",x"70",x"80",x"c1"),
   536 => (x"ff",x"05",x"8d",x"c1"),
   537 => (x"d0",x"ff",x"87",x"f0"),
   538 => (x"72",x"78",x"c4",x"48"),
   539 => (x"c5",x"c0",x"05",x"9a"),
   540 => (x"c0",x"48",x"c0",x"87"),
   541 => (x"1e",x"c1",x"87",x"e6"),
   542 => (x"49",x"f2",x"f6",x"c2"),
   543 => (x"87",x"dd",x"ff",x"fd"),
   544 => (x"9c",x"74",x"86",x"c4"),
   545 => (x"87",x"c3",x"fe",x"05"),
   546 => (x"c8",x"48",x"d0",x"ff"),
   547 => (x"d3",x"c1",x"78",x"c5"),
   548 => (x"c4",x"7b",x"c0",x"7b"),
   549 => (x"c0",x"48",x"c1",x"78"),
   550 => (x"48",x"c0",x"87",x"c2"),
   551 => (x"26",x"4d",x"26",x"26"),
   552 => (x"26",x"4b",x"26",x"4c"),
   553 => (x"4a",x"71",x"1e",x"4f"),
   554 => (x"c5",x"05",x"66",x"c4"),
   555 => (x"fb",x"49",x"72",x"87"),
   556 => (x"4f",x"26",x"87",x"ca"),
   557 => (x"e4",x"c2",x"1e",x"00"),
   558 => (x"c1",x"49",x"bf",x"c3"),
   559 => (x"c7",x"e4",x"c2",x"b9"),
   560 => (x"48",x"d4",x"ff",x"59"),
   561 => (x"ff",x"78",x"ff",x"c3"),
   562 => (x"e1",x"c8",x"48",x"d0"),
   563 => (x"48",x"d4",x"ff",x"78"),
   564 => (x"31",x"c4",x"78",x"c1"),
   565 => (x"d0",x"ff",x"78",x"71"),
   566 => (x"78",x"e0",x"c0",x"48"),
   567 => (x"c2",x"1e",x"4f",x"26"),
   568 => (x"c2",x"1e",x"f7",x"e3"),
   569 => (x"fd",x"49",x"f2",x"f6"),
   570 => (x"c4",x"87",x"f7",x"fb"),
   571 => (x"02",x"98",x"70",x"86"),
   572 => (x"c0",x"ff",x"87",x"c3"),
   573 => (x"31",x"4f",x"26",x"87"),
   574 => (x"5a",x"48",x"4b",x"35"),
   575 => (x"43",x"20",x"20",x"20"),
   576 => (x"00",x"00",x"47",x"46"),
   577 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

