
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c8",x"f7",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"c8",x"f7",x"c2"),
    14 => (x"48",x"c8",x"e4",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e1",x"e0"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"ff",x"1e",x"4f",x"26"),
    53 => (x"ff",x"c3",x"48",x"d4"),
    54 => (x"c4",x"51",x"68",x"78"),
    55 => (x"88",x"c1",x"48",x"66"),
    56 => (x"70",x"58",x"a6",x"c8"),
    57 => (x"87",x"eb",x"05",x"98"),
    58 => (x"73",x"1e",x"4f",x"26"),
    59 => (x"4b",x"d4",x"ff",x"1e"),
    60 => (x"6b",x"7b",x"ff",x"c3"),
    61 => (x"7b",x"ff",x"c3",x"4a"),
    62 => (x"32",x"c8",x"49",x"6b"),
    63 => (x"ff",x"c3",x"b1",x"72"),
    64 => (x"c8",x"4a",x"6b",x"7b"),
    65 => (x"c3",x"b2",x"71",x"31"),
    66 => (x"49",x"6b",x"7b",x"ff"),
    67 => (x"b1",x"72",x"32",x"c8"),
    68 => (x"87",x"c4",x"48",x"71"),
    69 => (x"4c",x"26",x"4d",x"26"),
    70 => (x"4f",x"26",x"4b",x"26"),
    71 => (x"5c",x"5b",x"5e",x"0e"),
    72 => (x"4a",x"71",x"0e",x"5d"),
    73 => (x"72",x"4c",x"d4",x"ff"),
    74 => (x"99",x"ff",x"c3",x"49"),
    75 => (x"e4",x"c2",x"7c",x"71"),
    76 => (x"c8",x"05",x"bf",x"c8"),
    77 => (x"48",x"66",x"d0",x"87"),
    78 => (x"a6",x"d4",x"30",x"c9"),
    79 => (x"49",x"66",x"d0",x"58"),
    80 => (x"ff",x"c3",x"29",x"d8"),
    81 => (x"d0",x"7c",x"71",x"99"),
    82 => (x"29",x"d0",x"49",x"66"),
    83 => (x"71",x"99",x"ff",x"c3"),
    84 => (x"49",x"66",x"d0",x"7c"),
    85 => (x"ff",x"c3",x"29",x"c8"),
    86 => (x"d0",x"7c",x"71",x"99"),
    87 => (x"ff",x"c3",x"49",x"66"),
    88 => (x"72",x"7c",x"71",x"99"),
    89 => (x"c3",x"29",x"d0",x"49"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"f0",x"c9",x"4b",x"6c"),
    92 => (x"ff",x"c3",x"4d",x"ff"),
    93 => (x"87",x"d0",x"05",x"ab"),
    94 => (x"6c",x"7c",x"ff",x"c3"),
    95 => (x"02",x"8d",x"c1",x"4b"),
    96 => (x"ff",x"c3",x"87",x"c6"),
    97 => (x"87",x"f0",x"02",x"ab"),
    98 => (x"c7",x"fe",x"48",x"73"),
    99 => (x"49",x"c0",x"1e",x"87"),
   100 => (x"c3",x"48",x"d4",x"ff"),
   101 => (x"81",x"c1",x"78",x"ff"),
   102 => (x"a9",x"b7",x"c8",x"c3"),
   103 => (x"26",x"87",x"f1",x"04"),
   104 => (x"1e",x"73",x"1e",x"4f"),
   105 => (x"f8",x"c4",x"87",x"e7"),
   106 => (x"1e",x"c0",x"4b",x"df"),
   107 => (x"c1",x"f0",x"ff",x"c0"),
   108 => (x"e7",x"fd",x"49",x"f7"),
   109 => (x"c1",x"86",x"c4",x"87"),
   110 => (x"ea",x"c0",x"05",x"a8"),
   111 => (x"48",x"d4",x"ff",x"87"),
   112 => (x"c1",x"78",x"ff",x"c3"),
   113 => (x"c0",x"c0",x"c0",x"c0"),
   114 => (x"e1",x"c0",x"1e",x"c0"),
   115 => (x"49",x"e9",x"c1",x"f0"),
   116 => (x"c4",x"87",x"c9",x"fd"),
   117 => (x"05",x"98",x"70",x"86"),
   118 => (x"d4",x"ff",x"87",x"ca"),
   119 => (x"78",x"ff",x"c3",x"48"),
   120 => (x"87",x"cb",x"48",x"c1"),
   121 => (x"c1",x"87",x"e6",x"fe"),
   122 => (x"fd",x"fe",x"05",x"8b"),
   123 => (x"fc",x"48",x"c0",x"87"),
   124 => (x"73",x"1e",x"87",x"e6"),
   125 => (x"48",x"d4",x"ff",x"1e"),
   126 => (x"d3",x"78",x"ff",x"c3"),
   127 => (x"c0",x"1e",x"c0",x"4b"),
   128 => (x"c1",x"c1",x"f0",x"ff"),
   129 => (x"87",x"d4",x"fc",x"49"),
   130 => (x"98",x"70",x"86",x"c4"),
   131 => (x"ff",x"87",x"ca",x"05"),
   132 => (x"ff",x"c3",x"48",x"d4"),
   133 => (x"cb",x"48",x"c1",x"78"),
   134 => (x"87",x"f1",x"fd",x"87"),
   135 => (x"ff",x"05",x"8b",x"c1"),
   136 => (x"48",x"c0",x"87",x"db"),
   137 => (x"0e",x"87",x"f1",x"fb"),
   138 => (x"0e",x"5c",x"5b",x"5e"),
   139 => (x"fd",x"4c",x"d4",x"ff"),
   140 => (x"ea",x"c6",x"87",x"db"),
   141 => (x"f0",x"e1",x"c0",x"1e"),
   142 => (x"fb",x"49",x"c8",x"c1"),
   143 => (x"86",x"c4",x"87",x"de"),
   144 => (x"c8",x"02",x"a8",x"c1"),
   145 => (x"87",x"ea",x"fe",x"87"),
   146 => (x"e2",x"c1",x"48",x"c0"),
   147 => (x"87",x"da",x"fa",x"87"),
   148 => (x"ff",x"cf",x"49",x"70"),
   149 => (x"ea",x"c6",x"99",x"ff"),
   150 => (x"87",x"c8",x"02",x"a9"),
   151 => (x"c0",x"87",x"d3",x"fe"),
   152 => (x"87",x"cb",x"c1",x"48"),
   153 => (x"c0",x"7c",x"ff",x"c3"),
   154 => (x"f4",x"fc",x"4b",x"f1"),
   155 => (x"02",x"98",x"70",x"87"),
   156 => (x"c0",x"87",x"eb",x"c0"),
   157 => (x"f0",x"ff",x"c0",x"1e"),
   158 => (x"fa",x"49",x"fa",x"c1"),
   159 => (x"86",x"c4",x"87",x"de"),
   160 => (x"d9",x"05",x"98",x"70"),
   161 => (x"7c",x"ff",x"c3",x"87"),
   162 => (x"ff",x"c3",x"49",x"6c"),
   163 => (x"7c",x"7c",x"7c",x"7c"),
   164 => (x"02",x"99",x"c0",x"c1"),
   165 => (x"48",x"c1",x"87",x"c4"),
   166 => (x"48",x"c0",x"87",x"d5"),
   167 => (x"ab",x"c2",x"87",x"d1"),
   168 => (x"c0",x"87",x"c4",x"05"),
   169 => (x"c1",x"87",x"c8",x"48"),
   170 => (x"fd",x"fe",x"05",x"8b"),
   171 => (x"f9",x"48",x"c0",x"87"),
   172 => (x"73",x"1e",x"87",x"e4"),
   173 => (x"c8",x"e4",x"c2",x"1e"),
   174 => (x"c7",x"78",x"c1",x"48"),
   175 => (x"48",x"d0",x"ff",x"4b"),
   176 => (x"c8",x"fb",x"78",x"c2"),
   177 => (x"48",x"d0",x"ff",x"87"),
   178 => (x"1e",x"c0",x"78",x"c3"),
   179 => (x"c1",x"d0",x"e5",x"c0"),
   180 => (x"c7",x"f9",x"49",x"c0"),
   181 => (x"c1",x"86",x"c4",x"87"),
   182 => (x"87",x"c1",x"05",x"a8"),
   183 => (x"05",x"ab",x"c2",x"4b"),
   184 => (x"48",x"c0",x"87",x"c5"),
   185 => (x"c1",x"87",x"f9",x"c0"),
   186 => (x"d0",x"ff",x"05",x"8b"),
   187 => (x"87",x"f7",x"fc",x"87"),
   188 => (x"58",x"cc",x"e4",x"c2"),
   189 => (x"cd",x"05",x"98",x"70"),
   190 => (x"c0",x"1e",x"c1",x"87"),
   191 => (x"d0",x"c1",x"f0",x"ff"),
   192 => (x"87",x"d8",x"f8",x"49"),
   193 => (x"d4",x"ff",x"86",x"c4"),
   194 => (x"78",x"ff",x"c3",x"48"),
   195 => (x"c2",x"87",x"fe",x"c2"),
   196 => (x"ff",x"58",x"d0",x"e4"),
   197 => (x"78",x"c2",x"48",x"d0"),
   198 => (x"c3",x"48",x"d4",x"ff"),
   199 => (x"48",x"c1",x"78",x"ff"),
   200 => (x"1e",x"87",x"f5",x"f7"),
   201 => (x"ff",x"4a",x"d4",x"ff"),
   202 => (x"d1",x"c4",x"48",x"d0"),
   203 => (x"7a",x"ff",x"c3",x"78"),
   204 => (x"f8",x"05",x"89",x"c1"),
   205 => (x"1e",x"4f",x"26",x"87"),
   206 => (x"4b",x"71",x"1e",x"73"),
   207 => (x"df",x"cd",x"ee",x"c5"),
   208 => (x"48",x"d4",x"ff",x"4a"),
   209 => (x"68",x"78",x"ff",x"c3"),
   210 => (x"a8",x"fe",x"c3",x"48"),
   211 => (x"c1",x"87",x"c5",x"02"),
   212 => (x"87",x"ed",x"05",x"8a"),
   213 => (x"c5",x"05",x"9a",x"72"),
   214 => (x"c0",x"48",x"c0",x"87"),
   215 => (x"9b",x"73",x"87",x"ea"),
   216 => (x"c8",x"87",x"cc",x"02"),
   217 => (x"49",x"73",x"1e",x"66"),
   218 => (x"c4",x"87",x"e7",x"f5"),
   219 => (x"c8",x"87",x"c6",x"86"),
   220 => (x"ee",x"fe",x"49",x"66"),
   221 => (x"48",x"d4",x"ff",x"87"),
   222 => (x"78",x"78",x"ff",x"c3"),
   223 => (x"c5",x"05",x"9b",x"73"),
   224 => (x"48",x"d0",x"ff",x"87"),
   225 => (x"48",x"c1",x"78",x"d0"),
   226 => (x"1e",x"87",x"cd",x"f6"),
   227 => (x"4a",x"71",x"1e",x"73"),
   228 => (x"d4",x"ff",x"4b",x"c0"),
   229 => (x"78",x"ff",x"c3",x"48"),
   230 => (x"c4",x"48",x"d0",x"ff"),
   231 => (x"d4",x"ff",x"78",x"c3"),
   232 => (x"78",x"ff",x"c3",x"48"),
   233 => (x"ff",x"c0",x"1e",x"72"),
   234 => (x"49",x"d1",x"c1",x"f0"),
   235 => (x"c4",x"87",x"ed",x"f5"),
   236 => (x"05",x"98",x"70",x"86"),
   237 => (x"c0",x"c8",x"87",x"cd"),
   238 => (x"49",x"66",x"cc",x"1e"),
   239 => (x"c4",x"87",x"f8",x"fd"),
   240 => (x"ff",x"4b",x"70",x"86"),
   241 => (x"78",x"c2",x"48",x"d0"),
   242 => (x"cb",x"f5",x"48",x"73"),
   243 => (x"5b",x"5e",x"0e",x"87"),
   244 => (x"c0",x"0e",x"5d",x"5c"),
   245 => (x"f0",x"ff",x"c0",x"1e"),
   246 => (x"f4",x"49",x"c9",x"c1"),
   247 => (x"1e",x"d2",x"87",x"fe"),
   248 => (x"49",x"d0",x"e4",x"c2"),
   249 => (x"c8",x"87",x"d0",x"fd"),
   250 => (x"c1",x"4c",x"c0",x"86"),
   251 => (x"ac",x"b7",x"d2",x"84"),
   252 => (x"c2",x"87",x"f8",x"04"),
   253 => (x"bf",x"97",x"d0",x"e4"),
   254 => (x"99",x"c0",x"c3",x"49"),
   255 => (x"05",x"a9",x"c0",x"c1"),
   256 => (x"c2",x"87",x"e7",x"c0"),
   257 => (x"bf",x"97",x"d7",x"e4"),
   258 => (x"c2",x"31",x"d0",x"49"),
   259 => (x"bf",x"97",x"d8",x"e4"),
   260 => (x"72",x"32",x"c8",x"4a"),
   261 => (x"d9",x"e4",x"c2",x"b1"),
   262 => (x"b1",x"4a",x"bf",x"97"),
   263 => (x"ff",x"cf",x"4c",x"71"),
   264 => (x"c1",x"9c",x"ff",x"ff"),
   265 => (x"c1",x"34",x"ca",x"84"),
   266 => (x"e4",x"c2",x"87",x"e7"),
   267 => (x"49",x"bf",x"97",x"d9"),
   268 => (x"99",x"c6",x"31",x"c1"),
   269 => (x"97",x"da",x"e4",x"c2"),
   270 => (x"b7",x"c7",x"4a",x"bf"),
   271 => (x"c2",x"b1",x"72",x"2a"),
   272 => (x"bf",x"97",x"d5",x"e4"),
   273 => (x"9d",x"cf",x"4d",x"4a"),
   274 => (x"97",x"d6",x"e4",x"c2"),
   275 => (x"9a",x"c3",x"4a",x"bf"),
   276 => (x"e4",x"c2",x"32",x"ca"),
   277 => (x"4b",x"bf",x"97",x"d7"),
   278 => (x"b2",x"73",x"33",x"c2"),
   279 => (x"97",x"d8",x"e4",x"c2"),
   280 => (x"c0",x"c3",x"4b",x"bf"),
   281 => (x"2b",x"b7",x"c6",x"9b"),
   282 => (x"81",x"c2",x"b2",x"73"),
   283 => (x"30",x"71",x"48",x"c1"),
   284 => (x"48",x"c1",x"49",x"70"),
   285 => (x"4d",x"70",x"30",x"75"),
   286 => (x"84",x"c1",x"4c",x"72"),
   287 => (x"c0",x"c8",x"94",x"71"),
   288 => (x"cc",x"06",x"ad",x"b7"),
   289 => (x"b7",x"34",x"c1",x"87"),
   290 => (x"b7",x"c0",x"c8",x"2d"),
   291 => (x"f4",x"ff",x"01",x"ad"),
   292 => (x"f1",x"48",x"74",x"87"),
   293 => (x"5e",x"0e",x"87",x"fe"),
   294 => (x"0e",x"5d",x"5c",x"5b"),
   295 => (x"ec",x"c2",x"86",x"f8"),
   296 => (x"78",x"c0",x"48",x"f6"),
   297 => (x"1e",x"ee",x"e4",x"c2"),
   298 => (x"de",x"fb",x"49",x"c0"),
   299 => (x"70",x"86",x"c4",x"87"),
   300 => (x"87",x"c5",x"05",x"98"),
   301 => (x"ce",x"c9",x"48",x"c0"),
   302 => (x"c1",x"4d",x"c0",x"87"),
   303 => (x"ca",x"f5",x"c0",x"7e"),
   304 => (x"e5",x"c2",x"49",x"bf"),
   305 => (x"c8",x"71",x"4a",x"e4"),
   306 => (x"87",x"de",x"ee",x"4b"),
   307 => (x"c2",x"05",x"98",x"70"),
   308 => (x"c0",x"7e",x"c0",x"87"),
   309 => (x"49",x"bf",x"c6",x"f5"),
   310 => (x"4a",x"c0",x"e6",x"c2"),
   311 => (x"ee",x"4b",x"c8",x"71"),
   312 => (x"98",x"70",x"87",x"c8"),
   313 => (x"c0",x"87",x"c2",x"05"),
   314 => (x"c0",x"02",x"6e",x"7e"),
   315 => (x"eb",x"c2",x"87",x"fd"),
   316 => (x"c2",x"4d",x"bf",x"f4"),
   317 => (x"bf",x"9f",x"ec",x"ec"),
   318 => (x"d6",x"c5",x"48",x"7e"),
   319 => (x"c7",x"05",x"a8",x"ea"),
   320 => (x"f4",x"eb",x"c2",x"87"),
   321 => (x"87",x"ce",x"4d",x"bf"),
   322 => (x"e9",x"ca",x"48",x"6e"),
   323 => (x"c5",x"02",x"a8",x"d5"),
   324 => (x"c7",x"48",x"c0",x"87"),
   325 => (x"e4",x"c2",x"87",x"f1"),
   326 => (x"49",x"75",x"1e",x"ee"),
   327 => (x"c4",x"87",x"ec",x"f9"),
   328 => (x"05",x"98",x"70",x"86"),
   329 => (x"48",x"c0",x"87",x"c5"),
   330 => (x"c0",x"87",x"dc",x"c7"),
   331 => (x"49",x"bf",x"c6",x"f5"),
   332 => (x"4a",x"c0",x"e6",x"c2"),
   333 => (x"ec",x"4b",x"c8",x"71"),
   334 => (x"98",x"70",x"87",x"f0"),
   335 => (x"c2",x"87",x"c8",x"05"),
   336 => (x"c1",x"48",x"f6",x"ec"),
   337 => (x"c0",x"87",x"da",x"78"),
   338 => (x"49",x"bf",x"ca",x"f5"),
   339 => (x"4a",x"e4",x"e5",x"c2"),
   340 => (x"ec",x"4b",x"c8",x"71"),
   341 => (x"98",x"70",x"87",x"d4"),
   342 => (x"87",x"c5",x"c0",x"02"),
   343 => (x"e6",x"c6",x"48",x"c0"),
   344 => (x"ec",x"ec",x"c2",x"87"),
   345 => (x"c1",x"49",x"bf",x"97"),
   346 => (x"c0",x"05",x"a9",x"d5"),
   347 => (x"ec",x"c2",x"87",x"cd"),
   348 => (x"49",x"bf",x"97",x"ed"),
   349 => (x"02",x"a9",x"ea",x"c2"),
   350 => (x"c0",x"87",x"c5",x"c0"),
   351 => (x"87",x"c7",x"c6",x"48"),
   352 => (x"97",x"ee",x"e4",x"c2"),
   353 => (x"c3",x"48",x"7e",x"bf"),
   354 => (x"c0",x"02",x"a8",x"e9"),
   355 => (x"48",x"6e",x"87",x"ce"),
   356 => (x"02",x"a8",x"eb",x"c3"),
   357 => (x"c0",x"87",x"c5",x"c0"),
   358 => (x"87",x"eb",x"c5",x"48"),
   359 => (x"97",x"f9",x"e4",x"c2"),
   360 => (x"05",x"99",x"49",x"bf"),
   361 => (x"c2",x"87",x"cc",x"c0"),
   362 => (x"bf",x"97",x"fa",x"e4"),
   363 => (x"02",x"a9",x"c2",x"49"),
   364 => (x"c0",x"87",x"c5",x"c0"),
   365 => (x"87",x"cf",x"c5",x"48"),
   366 => (x"97",x"fb",x"e4",x"c2"),
   367 => (x"ec",x"c2",x"48",x"bf"),
   368 => (x"4c",x"70",x"58",x"f2"),
   369 => (x"c2",x"88",x"c1",x"48"),
   370 => (x"c2",x"58",x"f6",x"ec"),
   371 => (x"bf",x"97",x"fc",x"e4"),
   372 => (x"c2",x"81",x"75",x"49"),
   373 => (x"bf",x"97",x"fd",x"e4"),
   374 => (x"72",x"32",x"c8",x"4a"),
   375 => (x"f1",x"c2",x"7e",x"a1"),
   376 => (x"78",x"6e",x"48",x"c3"),
   377 => (x"97",x"fe",x"e4",x"c2"),
   378 => (x"a6",x"c8",x"48",x"bf"),
   379 => (x"f6",x"ec",x"c2",x"58"),
   380 => (x"d4",x"c2",x"02",x"bf"),
   381 => (x"c6",x"f5",x"c0",x"87"),
   382 => (x"e6",x"c2",x"49",x"bf"),
   383 => (x"c8",x"71",x"4a",x"c0"),
   384 => (x"87",x"e6",x"e9",x"4b"),
   385 => (x"c0",x"02",x"98",x"70"),
   386 => (x"48",x"c0",x"87",x"c5"),
   387 => (x"c2",x"87",x"f8",x"c3"),
   388 => (x"4c",x"bf",x"ee",x"ec"),
   389 => (x"5c",x"d7",x"f1",x"c2"),
   390 => (x"97",x"d3",x"e5",x"c2"),
   391 => (x"31",x"c8",x"49",x"bf"),
   392 => (x"97",x"d2",x"e5",x"c2"),
   393 => (x"49",x"a1",x"4a",x"bf"),
   394 => (x"97",x"d4",x"e5",x"c2"),
   395 => (x"32",x"d0",x"4a",x"bf"),
   396 => (x"c2",x"49",x"a1",x"72"),
   397 => (x"bf",x"97",x"d5",x"e5"),
   398 => (x"72",x"32",x"d8",x"4a"),
   399 => (x"66",x"c4",x"49",x"a1"),
   400 => (x"c3",x"f1",x"c2",x"91"),
   401 => (x"f1",x"c2",x"81",x"bf"),
   402 => (x"e5",x"c2",x"59",x"cb"),
   403 => (x"4a",x"bf",x"97",x"db"),
   404 => (x"e5",x"c2",x"32",x"c8"),
   405 => (x"4b",x"bf",x"97",x"da"),
   406 => (x"e5",x"c2",x"4a",x"a2"),
   407 => (x"4b",x"bf",x"97",x"dc"),
   408 => (x"a2",x"73",x"33",x"d0"),
   409 => (x"dd",x"e5",x"c2",x"4a"),
   410 => (x"cf",x"4b",x"bf",x"97"),
   411 => (x"73",x"33",x"d8",x"9b"),
   412 => (x"f1",x"c2",x"4a",x"a2"),
   413 => (x"f1",x"c2",x"5a",x"cf"),
   414 => (x"c2",x"4a",x"bf",x"cb"),
   415 => (x"c2",x"92",x"74",x"8a"),
   416 => (x"72",x"48",x"cf",x"f1"),
   417 => (x"ca",x"c1",x"78",x"a1"),
   418 => (x"c0",x"e5",x"c2",x"87"),
   419 => (x"c8",x"49",x"bf",x"97"),
   420 => (x"ff",x"e4",x"c2",x"31"),
   421 => (x"a1",x"4a",x"bf",x"97"),
   422 => (x"fe",x"ec",x"c2",x"49"),
   423 => (x"fa",x"ec",x"c2",x"59"),
   424 => (x"31",x"c5",x"49",x"bf"),
   425 => (x"c9",x"81",x"ff",x"c7"),
   426 => (x"d7",x"f1",x"c2",x"29"),
   427 => (x"c5",x"e5",x"c2",x"59"),
   428 => (x"c8",x"4a",x"bf",x"97"),
   429 => (x"c4",x"e5",x"c2",x"32"),
   430 => (x"a2",x"4b",x"bf",x"97"),
   431 => (x"92",x"66",x"c4",x"4a"),
   432 => (x"f1",x"c2",x"82",x"6e"),
   433 => (x"f1",x"c2",x"5a",x"d3"),
   434 => (x"78",x"c0",x"48",x"cb"),
   435 => (x"48",x"c7",x"f1",x"c2"),
   436 => (x"c2",x"78",x"a1",x"72"),
   437 => (x"c2",x"48",x"d7",x"f1"),
   438 => (x"78",x"bf",x"cb",x"f1"),
   439 => (x"48",x"db",x"f1",x"c2"),
   440 => (x"bf",x"cf",x"f1",x"c2"),
   441 => (x"f6",x"ec",x"c2",x"78"),
   442 => (x"c9",x"c0",x"02",x"bf"),
   443 => (x"c4",x"48",x"74",x"87"),
   444 => (x"c0",x"7e",x"70",x"30"),
   445 => (x"f1",x"c2",x"87",x"c9"),
   446 => (x"c4",x"48",x"bf",x"d3"),
   447 => (x"c2",x"7e",x"70",x"30"),
   448 => (x"6e",x"48",x"fa",x"ec"),
   449 => (x"f8",x"48",x"c1",x"78"),
   450 => (x"26",x"4d",x"26",x"8e"),
   451 => (x"26",x"4b",x"26",x"4c"),
   452 => (x"5b",x"5e",x"0e",x"4f"),
   453 => (x"71",x"0e",x"5d",x"5c"),
   454 => (x"f6",x"ec",x"c2",x"4a"),
   455 => (x"87",x"cb",x"02",x"bf"),
   456 => (x"2b",x"c7",x"4b",x"72"),
   457 => (x"ff",x"c1",x"4c",x"72"),
   458 => (x"72",x"87",x"c9",x"9c"),
   459 => (x"72",x"2b",x"c8",x"4b"),
   460 => (x"9c",x"ff",x"c3",x"4c"),
   461 => (x"bf",x"c3",x"f1",x"c2"),
   462 => (x"c2",x"f5",x"c0",x"83"),
   463 => (x"d9",x"02",x"ab",x"bf"),
   464 => (x"c6",x"f5",x"c0",x"87"),
   465 => (x"ee",x"e4",x"c2",x"5b"),
   466 => (x"f0",x"49",x"73",x"1e"),
   467 => (x"86",x"c4",x"87",x"fd"),
   468 => (x"c5",x"05",x"98",x"70"),
   469 => (x"c0",x"48",x"c0",x"87"),
   470 => (x"ec",x"c2",x"87",x"e6"),
   471 => (x"d2",x"02",x"bf",x"f6"),
   472 => (x"c4",x"49",x"74",x"87"),
   473 => (x"ee",x"e4",x"c2",x"91"),
   474 => (x"cf",x"4d",x"69",x"81"),
   475 => (x"ff",x"ff",x"ff",x"ff"),
   476 => (x"74",x"87",x"cb",x"9d"),
   477 => (x"c2",x"91",x"c2",x"49"),
   478 => (x"9f",x"81",x"ee",x"e4"),
   479 => (x"48",x"75",x"4d",x"69"),
   480 => (x"0e",x"87",x"c6",x"fe"),
   481 => (x"5d",x"5c",x"5b",x"5e"),
   482 => (x"4d",x"71",x"1e",x"0e"),
   483 => (x"49",x"c1",x"1e",x"c0"),
   484 => (x"c4",x"87",x"d7",x"cf"),
   485 => (x"9c",x"4c",x"70",x"86"),
   486 => (x"87",x"c0",x"c1",x"02"),
   487 => (x"4a",x"fe",x"ec",x"c2"),
   488 => (x"ea",x"e2",x"49",x"75"),
   489 => (x"02",x"98",x"70",x"87"),
   490 => (x"74",x"87",x"f1",x"c0"),
   491 => (x"cb",x"49",x"75",x"4a"),
   492 => (x"87",x"d0",x"e3",x"4b"),
   493 => (x"c0",x"02",x"98",x"70"),
   494 => (x"1e",x"c0",x"87",x"e2"),
   495 => (x"c7",x"02",x"9c",x"74"),
   496 => (x"48",x"a6",x"c4",x"87"),
   497 => (x"87",x"c5",x"78",x"c0"),
   498 => (x"c1",x"48",x"a6",x"c4"),
   499 => (x"49",x"66",x"c4",x"78"),
   500 => (x"c4",x"87",x"d7",x"ce"),
   501 => (x"9c",x"4c",x"70",x"86"),
   502 => (x"87",x"c0",x"ff",x"05"),
   503 => (x"fc",x"26",x"48",x"74"),
   504 => (x"5e",x"0e",x"87",x"e7"),
   505 => (x"0e",x"5d",x"5c",x"5b"),
   506 => (x"9b",x"4b",x"71",x"1e"),
   507 => (x"c0",x"87",x"c5",x"05"),
   508 => (x"87",x"e5",x"c1",x"48"),
   509 => (x"c0",x"4d",x"a3",x"c8"),
   510 => (x"02",x"66",x"d4",x"7d"),
   511 => (x"66",x"d4",x"87",x"c7"),
   512 => (x"c5",x"05",x"bf",x"97"),
   513 => (x"c1",x"48",x"c0",x"87"),
   514 => (x"66",x"d4",x"87",x"cf"),
   515 => (x"87",x"f3",x"fd",x"49"),
   516 => (x"02",x"9c",x"4c",x"70"),
   517 => (x"dc",x"87",x"c0",x"c1"),
   518 => (x"7d",x"69",x"49",x"a4"),
   519 => (x"c4",x"49",x"a4",x"da"),
   520 => (x"69",x"9f",x"4a",x"a3"),
   521 => (x"f6",x"ec",x"c2",x"7a"),
   522 => (x"87",x"d2",x"02",x"bf"),
   523 => (x"9f",x"49",x"a4",x"d4"),
   524 => (x"ff",x"c0",x"49",x"69"),
   525 => (x"48",x"71",x"99",x"ff"),
   526 => (x"7e",x"70",x"30",x"d0"),
   527 => (x"7e",x"c0",x"87",x"c2"),
   528 => (x"6a",x"48",x"49",x"6e"),
   529 => (x"c0",x"7a",x"70",x"80"),
   530 => (x"49",x"a3",x"cc",x"7b"),
   531 => (x"a3",x"d0",x"79",x"6a"),
   532 => (x"74",x"79",x"c0",x"49"),
   533 => (x"c0",x"87",x"c2",x"48"),
   534 => (x"ec",x"fa",x"26",x"48"),
   535 => (x"5b",x"5e",x"0e",x"87"),
   536 => (x"71",x"0e",x"5d",x"5c"),
   537 => (x"c2",x"f5",x"c0",x"4c"),
   538 => (x"74",x"78",x"ff",x"48"),
   539 => (x"ca",x"c1",x"02",x"9c"),
   540 => (x"49",x"a4",x"c8",x"87"),
   541 => (x"c2",x"c1",x"02",x"69"),
   542 => (x"4a",x"66",x"d0",x"87"),
   543 => (x"d4",x"82",x"49",x"6c"),
   544 => (x"66",x"d0",x"5a",x"a6"),
   545 => (x"ec",x"c2",x"b9",x"4d"),
   546 => (x"ff",x"4a",x"bf",x"f2"),
   547 => (x"71",x"99",x"72",x"ba"),
   548 => (x"e4",x"c0",x"02",x"99"),
   549 => (x"4b",x"a4",x"c4",x"87"),
   550 => (x"f4",x"f9",x"49",x"6b"),
   551 => (x"c2",x"7b",x"70",x"87"),
   552 => (x"49",x"bf",x"ee",x"ec"),
   553 => (x"7c",x"71",x"81",x"6c"),
   554 => (x"ec",x"c2",x"b9",x"75"),
   555 => (x"ff",x"4a",x"bf",x"f2"),
   556 => (x"71",x"99",x"72",x"ba"),
   557 => (x"dc",x"ff",x"05",x"99"),
   558 => (x"f9",x"7c",x"75",x"87"),
   559 => (x"73",x"1e",x"87",x"cb"),
   560 => (x"9b",x"4b",x"71",x"1e"),
   561 => (x"c8",x"87",x"c7",x"02"),
   562 => (x"05",x"69",x"49",x"a3"),
   563 => (x"48",x"c0",x"87",x"c5"),
   564 => (x"c2",x"87",x"eb",x"c0"),
   565 => (x"4a",x"bf",x"c7",x"f1"),
   566 => (x"69",x"49",x"a3",x"c4"),
   567 => (x"c2",x"89",x"c2",x"49"),
   568 => (x"91",x"bf",x"ee",x"ec"),
   569 => (x"c2",x"4a",x"a2",x"71"),
   570 => (x"49",x"bf",x"f2",x"ec"),
   571 => (x"a2",x"71",x"99",x"6b"),
   572 => (x"1e",x"66",x"c8",x"4a"),
   573 => (x"d2",x"ea",x"49",x"72"),
   574 => (x"70",x"86",x"c4",x"87"),
   575 => (x"cc",x"f8",x"48",x"49"),
   576 => (x"5b",x"5e",x"0e",x"87"),
   577 => (x"1e",x"0e",x"5d",x"5c"),
   578 => (x"66",x"d4",x"4b",x"71"),
   579 => (x"73",x"2c",x"c9",x"4c"),
   580 => (x"cf",x"c1",x"02",x"9b"),
   581 => (x"49",x"a3",x"c8",x"87"),
   582 => (x"c7",x"c1",x"02",x"69"),
   583 => (x"4d",x"a3",x"d0",x"87"),
   584 => (x"c2",x"7d",x"66",x"d4"),
   585 => (x"49",x"bf",x"f2",x"ec"),
   586 => (x"4a",x"6b",x"b9",x"ff"),
   587 => (x"ac",x"71",x"7e",x"99"),
   588 => (x"c0",x"87",x"cd",x"03"),
   589 => (x"a3",x"cc",x"7d",x"7b"),
   590 => (x"49",x"a3",x"c4",x"4a"),
   591 => (x"87",x"c2",x"79",x"6a"),
   592 => (x"9c",x"74",x"8c",x"72"),
   593 => (x"49",x"87",x"dd",x"02"),
   594 => (x"fc",x"49",x"73",x"1e"),
   595 => (x"86",x"c4",x"87",x"cf"),
   596 => (x"c7",x"49",x"66",x"d4"),
   597 => (x"cb",x"02",x"99",x"ff"),
   598 => (x"ee",x"e4",x"c2",x"87"),
   599 => (x"fd",x"49",x"73",x"1e"),
   600 => (x"86",x"c4",x"87",x"dc"),
   601 => (x"87",x"e1",x"f6",x"26"),
   602 => (x"5c",x"5b",x"5e",x"0e"),
   603 => (x"86",x"f0",x"0e",x"5d"),
   604 => (x"c0",x"59",x"a6",x"d0"),
   605 => (x"cc",x"4b",x"66",x"e4"),
   606 => (x"87",x"ca",x"02",x"66"),
   607 => (x"70",x"80",x"c8",x"48"),
   608 => (x"05",x"bf",x"6e",x"7e"),
   609 => (x"48",x"c0",x"87",x"c5"),
   610 => (x"cc",x"87",x"ec",x"c3"),
   611 => (x"84",x"d0",x"4c",x"66"),
   612 => (x"a6",x"c4",x"49",x"73"),
   613 => (x"c4",x"78",x"6c",x"48"),
   614 => (x"80",x"c4",x"81",x"66"),
   615 => (x"c8",x"78",x"bf",x"6e"),
   616 => (x"c6",x"06",x"a9",x"66"),
   617 => (x"66",x"c4",x"49",x"87"),
   618 => (x"c0",x"4b",x"71",x"89"),
   619 => (x"c4",x"01",x"ab",x"b7"),
   620 => (x"c2",x"c3",x"48",x"87"),
   621 => (x"48",x"66",x"c4",x"87"),
   622 => (x"70",x"98",x"ff",x"c7"),
   623 => (x"c1",x"02",x"6e",x"7e"),
   624 => (x"c0",x"c8",x"87",x"c9"),
   625 => (x"71",x"89",x"6e",x"49"),
   626 => (x"ee",x"e4",x"c2",x"4a"),
   627 => (x"73",x"85",x"6e",x"4d"),
   628 => (x"c1",x"06",x"aa",x"b7"),
   629 => (x"49",x"72",x"4a",x"87"),
   630 => (x"80",x"66",x"c4",x"48"),
   631 => (x"8b",x"72",x"7c",x"70"),
   632 => (x"71",x"8a",x"c1",x"49"),
   633 => (x"87",x"d9",x"02",x"99"),
   634 => (x"48",x"66",x"e0",x"c0"),
   635 => (x"e0",x"c0",x"50",x"15"),
   636 => (x"80",x"c1",x"48",x"66"),
   637 => (x"58",x"a6",x"e4",x"c0"),
   638 => (x"8a",x"c1",x"49",x"72"),
   639 => (x"e7",x"05",x"99",x"71"),
   640 => (x"d0",x"1e",x"c1",x"87"),
   641 => (x"d4",x"f9",x"49",x"66"),
   642 => (x"c0",x"86",x"c4",x"87"),
   643 => (x"c1",x"06",x"ab",x"b7"),
   644 => (x"e0",x"c0",x"87",x"e3"),
   645 => (x"ff",x"c7",x"4d",x"66"),
   646 => (x"c0",x"06",x"ab",x"b7"),
   647 => (x"1e",x"75",x"87",x"e2"),
   648 => (x"fa",x"49",x"66",x"d0"),
   649 => (x"c0",x"c8",x"87",x"d8"),
   650 => (x"c8",x"48",x"6c",x"85"),
   651 => (x"7c",x"70",x"80",x"c0"),
   652 => (x"c1",x"8b",x"c0",x"c8"),
   653 => (x"49",x"66",x"d4",x"1e"),
   654 => (x"c8",x"87",x"e2",x"f8"),
   655 => (x"87",x"ee",x"c0",x"86"),
   656 => (x"1e",x"ee",x"e4",x"c2"),
   657 => (x"f9",x"49",x"66",x"d0"),
   658 => (x"86",x"c4",x"87",x"f4"),
   659 => (x"4a",x"ee",x"e4",x"c2"),
   660 => (x"6c",x"48",x"49",x"73"),
   661 => (x"73",x"7c",x"70",x"80"),
   662 => (x"71",x"8b",x"c1",x"49"),
   663 => (x"87",x"ce",x"02",x"99"),
   664 => (x"c1",x"7d",x"97",x"12"),
   665 => (x"c1",x"49",x"73",x"85"),
   666 => (x"05",x"99",x"71",x"8b"),
   667 => (x"b7",x"c0",x"87",x"f2"),
   668 => (x"e1",x"fe",x"01",x"ab"),
   669 => (x"f0",x"48",x"c1",x"87"),
   670 => (x"87",x"cd",x"f2",x"8e"),
   671 => (x"5c",x"5b",x"5e",x"0e"),
   672 => (x"4b",x"71",x"0e",x"5d"),
   673 => (x"87",x"c7",x"02",x"9b"),
   674 => (x"6d",x"4d",x"a3",x"c8"),
   675 => (x"ff",x"87",x"c5",x"05"),
   676 => (x"87",x"fd",x"c0",x"48"),
   677 => (x"6c",x"4c",x"a3",x"d0"),
   678 => (x"99",x"ff",x"c7",x"49"),
   679 => (x"6c",x"87",x"d8",x"05"),
   680 => (x"c1",x"87",x"c9",x"02"),
   681 => (x"f6",x"49",x"73",x"1e"),
   682 => (x"86",x"c4",x"87",x"f3"),
   683 => (x"1e",x"ee",x"e4",x"c2"),
   684 => (x"c9",x"f8",x"49",x"73"),
   685 => (x"6c",x"86",x"c4",x"87"),
   686 => (x"04",x"aa",x"6d",x"4a"),
   687 => (x"48",x"ff",x"87",x"c4"),
   688 => (x"a2",x"c1",x"87",x"cf"),
   689 => (x"c7",x"49",x"72",x"7c"),
   690 => (x"e4",x"c2",x"99",x"ff"),
   691 => (x"69",x"97",x"81",x"ee"),
   692 => (x"87",x"f5",x"f0",x"48"),
   693 => (x"71",x"1e",x"73",x"1e"),
   694 => (x"c0",x"02",x"9b",x"4b"),
   695 => (x"f1",x"c2",x"87",x"e4"),
   696 => (x"4a",x"73",x"5b",x"db"),
   697 => (x"ec",x"c2",x"8a",x"c2"),
   698 => (x"92",x"49",x"bf",x"ee"),
   699 => (x"bf",x"c7",x"f1",x"c2"),
   700 => (x"c2",x"80",x"72",x"48"),
   701 => (x"71",x"58",x"df",x"f1"),
   702 => (x"c2",x"30",x"c4",x"48"),
   703 => (x"c0",x"58",x"fe",x"ec"),
   704 => (x"f1",x"c2",x"87",x"ed"),
   705 => (x"f1",x"c2",x"48",x"d7"),
   706 => (x"c2",x"78",x"bf",x"cb"),
   707 => (x"c2",x"48",x"db",x"f1"),
   708 => (x"78",x"bf",x"cf",x"f1"),
   709 => (x"bf",x"f6",x"ec",x"c2"),
   710 => (x"c2",x"87",x"c9",x"02"),
   711 => (x"49",x"bf",x"ee",x"ec"),
   712 => (x"87",x"c7",x"31",x"c4"),
   713 => (x"bf",x"d3",x"f1",x"c2"),
   714 => (x"c2",x"31",x"c4",x"49"),
   715 => (x"ef",x"59",x"fe",x"ec"),
   716 => (x"5e",x"0e",x"87",x"db"),
   717 => (x"71",x"0e",x"5c",x"5b"),
   718 => (x"72",x"4b",x"c0",x"4a"),
   719 => (x"e1",x"c0",x"02",x"9a"),
   720 => (x"49",x"a2",x"da",x"87"),
   721 => (x"c2",x"4b",x"69",x"9f"),
   722 => (x"02",x"bf",x"f6",x"ec"),
   723 => (x"a2",x"d4",x"87",x"cf"),
   724 => (x"49",x"69",x"9f",x"49"),
   725 => (x"ff",x"ff",x"c0",x"4c"),
   726 => (x"c2",x"34",x"d0",x"9c"),
   727 => (x"74",x"4c",x"c0",x"87"),
   728 => (x"49",x"73",x"b3",x"49"),
   729 => (x"ee",x"87",x"ed",x"fd"),
   730 => (x"5e",x"0e",x"87",x"e1"),
   731 => (x"0e",x"5d",x"5c",x"5b"),
   732 => (x"4a",x"71",x"86",x"f4"),
   733 => (x"9a",x"72",x"7e",x"c0"),
   734 => (x"c2",x"87",x"d8",x"02"),
   735 => (x"c0",x"48",x"ea",x"e4"),
   736 => (x"e2",x"e4",x"c2",x"78"),
   737 => (x"db",x"f1",x"c2",x"48"),
   738 => (x"e4",x"c2",x"78",x"bf"),
   739 => (x"f1",x"c2",x"48",x"e6"),
   740 => (x"c2",x"78",x"bf",x"d7"),
   741 => (x"c0",x"48",x"cb",x"ed"),
   742 => (x"fa",x"ec",x"c2",x"50"),
   743 => (x"e4",x"c2",x"49",x"bf"),
   744 => (x"71",x"4a",x"bf",x"ea"),
   745 => (x"c0",x"c4",x"03",x"aa"),
   746 => (x"cf",x"49",x"72",x"87"),
   747 => (x"e1",x"c0",x"05",x"99"),
   748 => (x"ee",x"e4",x"c2",x"87"),
   749 => (x"e2",x"e4",x"c2",x"1e"),
   750 => (x"e4",x"c2",x"49",x"bf"),
   751 => (x"a1",x"c1",x"48",x"e2"),
   752 => (x"df",x"ff",x"71",x"78"),
   753 => (x"86",x"c4",x"87",x"c5"),
   754 => (x"48",x"fe",x"f4",x"c0"),
   755 => (x"78",x"ee",x"e4",x"c2"),
   756 => (x"f4",x"c0",x"87",x"cc"),
   757 => (x"c0",x"48",x"bf",x"fe"),
   758 => (x"f5",x"c0",x"80",x"e0"),
   759 => (x"e4",x"c2",x"58",x"c2"),
   760 => (x"c1",x"48",x"bf",x"ea"),
   761 => (x"ee",x"e4",x"c2",x"80"),
   762 => (x"0d",x"3e",x"27",x"58"),
   763 => (x"97",x"bf",x"00",x"00"),
   764 => (x"02",x"9d",x"4d",x"bf"),
   765 => (x"c3",x"87",x"e2",x"c2"),
   766 => (x"c2",x"02",x"ad",x"e5"),
   767 => (x"f4",x"c0",x"87",x"db"),
   768 => (x"cb",x"4b",x"bf",x"fe"),
   769 => (x"4c",x"11",x"49",x"a3"),
   770 => (x"c1",x"05",x"ac",x"cf"),
   771 => (x"49",x"75",x"87",x"d2"),
   772 => (x"89",x"c1",x"99",x"df"),
   773 => (x"ec",x"c2",x"91",x"cd"),
   774 => (x"a3",x"c1",x"81",x"fe"),
   775 => (x"c3",x"51",x"12",x"4a"),
   776 => (x"51",x"12",x"4a",x"a3"),
   777 => (x"12",x"4a",x"a3",x"c5"),
   778 => (x"4a",x"a3",x"c7",x"51"),
   779 => (x"a3",x"c9",x"51",x"12"),
   780 => (x"ce",x"51",x"12",x"4a"),
   781 => (x"51",x"12",x"4a",x"a3"),
   782 => (x"12",x"4a",x"a3",x"d0"),
   783 => (x"4a",x"a3",x"d2",x"51"),
   784 => (x"a3",x"d4",x"51",x"12"),
   785 => (x"d6",x"51",x"12",x"4a"),
   786 => (x"51",x"12",x"4a",x"a3"),
   787 => (x"12",x"4a",x"a3",x"d8"),
   788 => (x"4a",x"a3",x"dc",x"51"),
   789 => (x"a3",x"de",x"51",x"12"),
   790 => (x"c1",x"51",x"12",x"4a"),
   791 => (x"87",x"f9",x"c0",x"7e"),
   792 => (x"99",x"c8",x"49",x"74"),
   793 => (x"87",x"ea",x"c0",x"05"),
   794 => (x"99",x"d0",x"49",x"74"),
   795 => (x"dc",x"87",x"d0",x"05"),
   796 => (x"ca",x"c0",x"02",x"66"),
   797 => (x"dc",x"49",x"73",x"87"),
   798 => (x"98",x"70",x"0f",x"66"),
   799 => (x"6e",x"87",x"d3",x"02"),
   800 => (x"87",x"c6",x"c0",x"05"),
   801 => (x"48",x"fe",x"ec",x"c2"),
   802 => (x"f4",x"c0",x"50",x"c0"),
   803 => (x"c2",x"48",x"bf",x"fe"),
   804 => (x"ed",x"c2",x"87",x"e7"),
   805 => (x"50",x"c0",x"48",x"cb"),
   806 => (x"fa",x"ec",x"c2",x"7e"),
   807 => (x"e4",x"c2",x"49",x"bf"),
   808 => (x"71",x"4a",x"bf",x"ea"),
   809 => (x"c0",x"fc",x"04",x"aa"),
   810 => (x"db",x"f1",x"c2",x"87"),
   811 => (x"c8",x"c0",x"05",x"bf"),
   812 => (x"f6",x"ec",x"c2",x"87"),
   813 => (x"fe",x"c1",x"02",x"bf"),
   814 => (x"c2",x"f5",x"c0",x"87"),
   815 => (x"c2",x"78",x"ff",x"48"),
   816 => (x"49",x"bf",x"e6",x"e4"),
   817 => (x"70",x"87",x"ca",x"e9"),
   818 => (x"ea",x"e4",x"c2",x"49"),
   819 => (x"48",x"a6",x"c4",x"59"),
   820 => (x"bf",x"e6",x"e4",x"c2"),
   821 => (x"f6",x"ec",x"c2",x"78"),
   822 => (x"d8",x"c0",x"02",x"bf"),
   823 => (x"49",x"66",x"c4",x"87"),
   824 => (x"ff",x"ff",x"ff",x"cf"),
   825 => (x"02",x"a9",x"99",x"f8"),
   826 => (x"c0",x"87",x"c5",x"c0"),
   827 => (x"87",x"e1",x"c0",x"4d"),
   828 => (x"dc",x"c0",x"4d",x"c1"),
   829 => (x"49",x"66",x"c4",x"87"),
   830 => (x"99",x"f8",x"ff",x"cf"),
   831 => (x"c8",x"c0",x"02",x"a9"),
   832 => (x"48",x"a6",x"c8",x"87"),
   833 => (x"c5",x"c0",x"78",x"c0"),
   834 => (x"48",x"a6",x"c8",x"87"),
   835 => (x"66",x"c8",x"78",x"c1"),
   836 => (x"05",x"9d",x"75",x"4d"),
   837 => (x"c4",x"87",x"e0",x"c0"),
   838 => (x"89",x"c2",x"49",x"66"),
   839 => (x"bf",x"ee",x"ec",x"c2"),
   840 => (x"f1",x"c2",x"91",x"4a"),
   841 => (x"c2",x"4a",x"bf",x"c7"),
   842 => (x"72",x"48",x"e2",x"e4"),
   843 => (x"e4",x"c2",x"78",x"a1"),
   844 => (x"78",x"c0",x"48",x"ea"),
   845 => (x"c0",x"87",x"e2",x"f9"),
   846 => (x"e7",x"8e",x"f4",x"48"),
   847 => (x"00",x"00",x"87",x"cb"),
   848 => (x"ff",x"ff",x"00",x"00"),
   849 => (x"0d",x"4e",x"ff",x"ff"),
   850 => (x"0d",x"57",x"00",x"00"),
   851 => (x"41",x"46",x"00",x"00"),
   852 => (x"20",x"32",x"33",x"54"),
   853 => (x"46",x"00",x"20",x"20"),
   854 => (x"36",x"31",x"54",x"41"),
   855 => (x"00",x"20",x"20",x"20"),
   856 => (x"e0",x"f1",x"c2",x"1e"),
   857 => (x"a8",x"dd",x"48",x"bf"),
   858 => (x"c0",x"87",x"c9",x"05"),
   859 => (x"70",x"87",x"d0",x"ff"),
   860 => (x"87",x"c8",x"4a",x"49"),
   861 => (x"c3",x"48",x"d4",x"ff"),
   862 => (x"4a",x"68",x"78",x"ff"),
   863 => (x"4f",x"26",x"48",x"72"),
   864 => (x"e0",x"f1",x"c2",x"1e"),
   865 => (x"a8",x"dd",x"48",x"bf"),
   866 => (x"c0",x"87",x"c6",x"05"),
   867 => (x"d9",x"87",x"dc",x"fe"),
   868 => (x"48",x"d4",x"ff",x"87"),
   869 => (x"ff",x"78",x"ff",x"c3"),
   870 => (x"e1",x"c8",x"48",x"d0"),
   871 => (x"48",x"d4",x"ff",x"78"),
   872 => (x"f1",x"c2",x"78",x"d4"),
   873 => (x"d4",x"ff",x"48",x"df"),
   874 => (x"4f",x"26",x"50",x"bf"),
   875 => (x"48",x"d0",x"ff",x"1e"),
   876 => (x"26",x"78",x"e0",x"c0"),
   877 => (x"e7",x"fe",x"1e",x"4f"),
   878 => (x"99",x"49",x"70",x"87"),
   879 => (x"c0",x"87",x"c6",x"02"),
   880 => (x"f1",x"05",x"a9",x"fb"),
   881 => (x"26",x"48",x"71",x"87"),
   882 => (x"5b",x"5e",x"0e",x"4f"),
   883 => (x"4b",x"71",x"0e",x"5c"),
   884 => (x"cb",x"fe",x"4c",x"c0"),
   885 => (x"99",x"49",x"70",x"87"),
   886 => (x"87",x"f9",x"c0",x"02"),
   887 => (x"02",x"a9",x"ec",x"c0"),
   888 => (x"c0",x"87",x"f2",x"c0"),
   889 => (x"c0",x"02",x"a9",x"fb"),
   890 => (x"66",x"cc",x"87",x"eb"),
   891 => (x"c7",x"03",x"ac",x"b7"),
   892 => (x"02",x"66",x"d0",x"87"),
   893 => (x"53",x"71",x"87",x"c2"),
   894 => (x"c2",x"02",x"99",x"71"),
   895 => (x"fd",x"84",x"c1",x"87"),
   896 => (x"49",x"70",x"87",x"de"),
   897 => (x"87",x"cd",x"02",x"99"),
   898 => (x"02",x"a9",x"ec",x"c0"),
   899 => (x"fb",x"c0",x"87",x"c7"),
   900 => (x"d5",x"ff",x"05",x"a9"),
   901 => (x"02",x"66",x"d0",x"87"),
   902 => (x"97",x"c0",x"87",x"c3"),
   903 => (x"a9",x"ec",x"c0",x"7b"),
   904 => (x"74",x"87",x"c4",x"05"),
   905 => (x"74",x"87",x"c5",x"4a"),
   906 => (x"8a",x"0a",x"c0",x"4a"),
   907 => (x"87",x"c2",x"48",x"72"),
   908 => (x"4c",x"26",x"4d",x"26"),
   909 => (x"4f",x"26",x"4b",x"26"),
   910 => (x"87",x"e4",x"fc",x"1e"),
   911 => (x"f0",x"c0",x"49",x"70"),
   912 => (x"ca",x"04",x"a9",x"b7"),
   913 => (x"b7",x"f9",x"c0",x"87"),
   914 => (x"87",x"c3",x"01",x"a9"),
   915 => (x"c1",x"89",x"f0",x"c0"),
   916 => (x"04",x"a9",x"b7",x"c1"),
   917 => (x"da",x"c1",x"87",x"ca"),
   918 => (x"c3",x"01",x"a9",x"b7"),
   919 => (x"89",x"f7",x"c0",x"87"),
   920 => (x"4f",x"26",x"48",x"71"),
   921 => (x"5c",x"5b",x"5e",x"0e"),
   922 => (x"ff",x"4a",x"71",x"0e"),
   923 => (x"49",x"72",x"4c",x"d4"),
   924 => (x"70",x"87",x"ea",x"c0"),
   925 => (x"c2",x"02",x"9b",x"4b"),
   926 => (x"ff",x"8b",x"c1",x"87"),
   927 => (x"c5",x"c8",x"48",x"d0"),
   928 => (x"7c",x"d5",x"c1",x"78"),
   929 => (x"31",x"c6",x"49",x"73"),
   930 => (x"97",x"f4",x"e2",x"c2"),
   931 => (x"71",x"48",x"4a",x"bf"),
   932 => (x"ff",x"7c",x"70",x"b0"),
   933 => (x"78",x"c4",x"48",x"d0"),
   934 => (x"d5",x"fe",x"48",x"73"),
   935 => (x"5b",x"5e",x"0e",x"87"),
   936 => (x"f4",x"0e",x"5d",x"5c"),
   937 => (x"c4",x"4c",x"71",x"86"),
   938 => (x"78",x"c0",x"48",x"a6"),
   939 => (x"6e",x"7e",x"a4",x"c8"),
   940 => (x"c1",x"49",x"bf",x"97"),
   941 => (x"dd",x"05",x"a9",x"c1"),
   942 => (x"49",x"a4",x"c9",x"87"),
   943 => (x"c1",x"49",x"69",x"97"),
   944 => (x"d1",x"05",x"a9",x"d2"),
   945 => (x"49",x"a4",x"ca",x"87"),
   946 => (x"c1",x"49",x"69",x"97"),
   947 => (x"c5",x"05",x"a9",x"c3"),
   948 => (x"c2",x"48",x"df",x"87"),
   949 => (x"e7",x"fa",x"87",x"e1"),
   950 => (x"c0",x"4b",x"c0",x"87"),
   951 => (x"bf",x"97",x"fc",x"fd"),
   952 => (x"04",x"a9",x"c0",x"49"),
   953 => (x"cc",x"fb",x"87",x"cf"),
   954 => (x"c0",x"83",x"c1",x"87"),
   955 => (x"bf",x"97",x"fc",x"fd"),
   956 => (x"f1",x"06",x"ab",x"49"),
   957 => (x"fc",x"fd",x"c0",x"87"),
   958 => (x"cf",x"02",x"bf",x"97"),
   959 => (x"87",x"e0",x"f9",x"87"),
   960 => (x"02",x"99",x"49",x"70"),
   961 => (x"ec",x"c0",x"87",x"c6"),
   962 => (x"87",x"f1",x"05",x"a9"),
   963 => (x"cf",x"f9",x"4b",x"c0"),
   964 => (x"f9",x"4d",x"70",x"87"),
   965 => (x"a6",x"cc",x"87",x"ca"),
   966 => (x"87",x"c4",x"f9",x"58"),
   967 => (x"83",x"c1",x"4a",x"70"),
   968 => (x"49",x"bf",x"97",x"6e"),
   969 => (x"87",x"c7",x"02",x"ad"),
   970 => (x"05",x"ad",x"ff",x"c0"),
   971 => (x"c9",x"87",x"ea",x"c0"),
   972 => (x"69",x"97",x"49",x"a4"),
   973 => (x"a9",x"66",x"c8",x"49"),
   974 => (x"48",x"87",x"c7",x"02"),
   975 => (x"05",x"a8",x"ff",x"c0"),
   976 => (x"a4",x"ca",x"87",x"d7"),
   977 => (x"49",x"69",x"97",x"49"),
   978 => (x"87",x"c6",x"02",x"aa"),
   979 => (x"05",x"aa",x"ff",x"c0"),
   980 => (x"a6",x"c4",x"87",x"c7"),
   981 => (x"d3",x"78",x"c1",x"48"),
   982 => (x"ad",x"ec",x"c0",x"87"),
   983 => (x"c0",x"87",x"c6",x"02"),
   984 => (x"c7",x"05",x"ad",x"fb"),
   985 => (x"c4",x"4b",x"c0",x"87"),
   986 => (x"78",x"c1",x"48",x"a6"),
   987 => (x"fe",x"02",x"66",x"c4"),
   988 => (x"f7",x"f8",x"87",x"dc"),
   989 => (x"f4",x"48",x"73",x"87"),
   990 => (x"87",x"f4",x"fa",x"8e"),
   991 => (x"5b",x"5e",x"0e",x"00"),
   992 => (x"1e",x"0e",x"5d",x"5c"),
   993 => (x"4c",x"c0",x"4b",x"71"),
   994 => (x"c0",x"04",x"ab",x"4d"),
   995 => (x"fa",x"c0",x"87",x"e8"),
   996 => (x"9d",x"75",x"1e",x"dd"),
   997 => (x"c0",x"87",x"c4",x"02"),
   998 => (x"c1",x"87",x"c2",x"4a"),
   999 => (x"ef",x"49",x"72",x"4a"),
  1000 => (x"86",x"c4",x"87",x"c8"),
  1001 => (x"84",x"c1",x"7e",x"70"),
  1002 => (x"87",x"c2",x"05",x"6e"),
  1003 => (x"85",x"c1",x"4c",x"73"),
  1004 => (x"ff",x"06",x"ac",x"73"),
  1005 => (x"48",x"6e",x"87",x"d8"),
  1006 => (x"26",x"4d",x"26",x"26"),
  1007 => (x"26",x"4b",x"26",x"4c"),
  1008 => (x"5b",x"5e",x"0e",x"4f"),
  1009 => (x"1e",x"0e",x"5d",x"5c"),
  1010 => (x"de",x"49",x"4c",x"71"),
  1011 => (x"f9",x"f1",x"c2",x"91"),
  1012 => (x"97",x"85",x"71",x"4d"),
  1013 => (x"dd",x"c1",x"02",x"6d"),
  1014 => (x"e4",x"f1",x"c2",x"87"),
  1015 => (x"82",x"74",x"4a",x"bf"),
  1016 => (x"d8",x"fe",x"49",x"72"),
  1017 => (x"6e",x"7e",x"70",x"87"),
  1018 => (x"87",x"f3",x"c0",x"02"),
  1019 => (x"4b",x"ec",x"f1",x"c2"),
  1020 => (x"49",x"cb",x"4a",x"6e"),
  1021 => (x"87",x"f0",x"c2",x"ff"),
  1022 => (x"93",x"cb",x"4b",x"74"),
  1023 => (x"83",x"d0",x"e2",x"c1"),
  1024 => (x"c0",x"c1",x"83",x"c4"),
  1025 => (x"49",x"74",x"7b",x"fa"),
  1026 => (x"87",x"fe",x"cd",x"c1"),
  1027 => (x"f1",x"c2",x"7b",x"75"),
  1028 => (x"49",x"bf",x"97",x"f8"),
  1029 => (x"ec",x"f1",x"c2",x"1e"),
  1030 => (x"c8",x"e2",x"c1",x"49"),
  1031 => (x"74",x"86",x"c4",x"87"),
  1032 => (x"e5",x"cd",x"c1",x"49"),
  1033 => (x"c1",x"49",x"c0",x"87"),
  1034 => (x"c2",x"87",x"c4",x"cf"),
  1035 => (x"c0",x"48",x"e0",x"f1"),
  1036 => (x"dd",x"49",x"c1",x"78"),
  1037 => (x"fd",x"26",x"87",x"cf"),
  1038 => (x"6f",x"4c",x"87",x"ff"),
  1039 => (x"6e",x"69",x"64",x"61"),
  1040 => (x"2e",x"2e",x"2e",x"67"),
  1041 => (x"5b",x"5e",x"0e",x"00"),
  1042 => (x"4b",x"71",x"0e",x"5c"),
  1043 => (x"e4",x"f1",x"c2",x"4a"),
  1044 => (x"49",x"72",x"82",x"bf"),
  1045 => (x"70",x"87",x"e6",x"fc"),
  1046 => (x"c4",x"02",x"9c",x"4c"),
  1047 => (x"d1",x"eb",x"49",x"87"),
  1048 => (x"e4",x"f1",x"c2",x"87"),
  1049 => (x"c1",x"78",x"c0",x"48"),
  1050 => (x"87",x"d9",x"dc",x"49"),
  1051 => (x"0e",x"87",x"cc",x"fd"),
  1052 => (x"5d",x"5c",x"5b",x"5e"),
  1053 => (x"c2",x"86",x"f4",x"0e"),
  1054 => (x"c0",x"4d",x"ee",x"e4"),
  1055 => (x"48",x"a6",x"c4",x"4c"),
  1056 => (x"f1",x"c2",x"78",x"c0"),
  1057 => (x"c0",x"49",x"bf",x"e4"),
  1058 => (x"c1",x"c1",x"06",x"a9"),
  1059 => (x"ee",x"e4",x"c2",x"87"),
  1060 => (x"c0",x"02",x"98",x"48"),
  1061 => (x"fa",x"c0",x"87",x"f8"),
  1062 => (x"66",x"c8",x"1e",x"dd"),
  1063 => (x"c4",x"87",x"c7",x"02"),
  1064 => (x"78",x"c0",x"48",x"a6"),
  1065 => (x"a6",x"c4",x"87",x"c5"),
  1066 => (x"c4",x"78",x"c1",x"48"),
  1067 => (x"f9",x"ea",x"49",x"66"),
  1068 => (x"70",x"86",x"c4",x"87"),
  1069 => (x"c4",x"84",x"c1",x"4d"),
  1070 => (x"80",x"c1",x"48",x"66"),
  1071 => (x"c2",x"58",x"a6",x"c8"),
  1072 => (x"49",x"bf",x"e4",x"f1"),
  1073 => (x"87",x"c6",x"03",x"ac"),
  1074 => (x"ff",x"05",x"9d",x"75"),
  1075 => (x"4c",x"c0",x"87",x"c8"),
  1076 => (x"c3",x"02",x"9d",x"75"),
  1077 => (x"fa",x"c0",x"87",x"e0"),
  1078 => (x"66",x"c8",x"1e",x"dd"),
  1079 => (x"cc",x"87",x"c7",x"02"),
  1080 => (x"78",x"c0",x"48",x"a6"),
  1081 => (x"a6",x"cc",x"87",x"c5"),
  1082 => (x"cc",x"78",x"c1",x"48"),
  1083 => (x"f9",x"e9",x"49",x"66"),
  1084 => (x"70",x"86",x"c4",x"87"),
  1085 => (x"c2",x"02",x"6e",x"7e"),
  1086 => (x"49",x"6e",x"87",x"e9"),
  1087 => (x"69",x"97",x"81",x"cb"),
  1088 => (x"02",x"99",x"d0",x"49"),
  1089 => (x"c1",x"87",x"d6",x"c1"),
  1090 => (x"74",x"4a",x"c5",x"c1"),
  1091 => (x"c1",x"91",x"cb",x"49"),
  1092 => (x"72",x"81",x"d0",x"e2"),
  1093 => (x"c3",x"81",x"c8",x"79"),
  1094 => (x"49",x"74",x"51",x"ff"),
  1095 => (x"f1",x"c2",x"91",x"de"),
  1096 => (x"85",x"71",x"4d",x"f9"),
  1097 => (x"7d",x"97",x"c1",x"c2"),
  1098 => (x"c0",x"49",x"a5",x"c1"),
  1099 => (x"ec",x"c2",x"51",x"e0"),
  1100 => (x"02",x"bf",x"97",x"fe"),
  1101 => (x"84",x"c1",x"87",x"d2"),
  1102 => (x"c2",x"4b",x"a5",x"c2"),
  1103 => (x"db",x"4a",x"fe",x"ec"),
  1104 => (x"e3",x"fd",x"fe",x"49"),
  1105 => (x"87",x"db",x"c1",x"87"),
  1106 => (x"c0",x"49",x"a5",x"cd"),
  1107 => (x"c2",x"84",x"c1",x"51"),
  1108 => (x"4a",x"6e",x"4b",x"a5"),
  1109 => (x"fd",x"fe",x"49",x"cb"),
  1110 => (x"c6",x"c1",x"87",x"ce"),
  1111 => (x"c1",x"ff",x"c0",x"87"),
  1112 => (x"cb",x"49",x"74",x"4a"),
  1113 => (x"d0",x"e2",x"c1",x"91"),
  1114 => (x"c2",x"79",x"72",x"81"),
  1115 => (x"bf",x"97",x"fe",x"ec"),
  1116 => (x"74",x"87",x"d8",x"02"),
  1117 => (x"c1",x"91",x"de",x"49"),
  1118 => (x"f9",x"f1",x"c2",x"84"),
  1119 => (x"c2",x"83",x"71",x"4b"),
  1120 => (x"dd",x"4a",x"fe",x"ec"),
  1121 => (x"df",x"fc",x"fe",x"49"),
  1122 => (x"74",x"87",x"d8",x"87"),
  1123 => (x"c2",x"93",x"de",x"4b"),
  1124 => (x"cb",x"83",x"f9",x"f1"),
  1125 => (x"51",x"c0",x"49",x"a3"),
  1126 => (x"6e",x"73",x"84",x"c1"),
  1127 => (x"fe",x"49",x"cb",x"4a"),
  1128 => (x"c4",x"87",x"c5",x"fc"),
  1129 => (x"80",x"c1",x"48",x"66"),
  1130 => (x"c7",x"58",x"a6",x"c8"),
  1131 => (x"c5",x"c0",x"03",x"ac"),
  1132 => (x"fc",x"05",x"6e",x"87"),
  1133 => (x"48",x"74",x"87",x"e0"),
  1134 => (x"fc",x"f7",x"8e",x"f4"),
  1135 => (x"1e",x"73",x"1e",x"87"),
  1136 => (x"cb",x"49",x"4b",x"71"),
  1137 => (x"d0",x"e2",x"c1",x"91"),
  1138 => (x"4a",x"a1",x"c8",x"81"),
  1139 => (x"48",x"f4",x"e2",x"c2"),
  1140 => (x"a1",x"c9",x"50",x"12"),
  1141 => (x"fc",x"fd",x"c0",x"4a"),
  1142 => (x"ca",x"50",x"12",x"48"),
  1143 => (x"f8",x"f1",x"c2",x"81"),
  1144 => (x"c2",x"50",x"11",x"48"),
  1145 => (x"bf",x"97",x"f8",x"f1"),
  1146 => (x"49",x"c0",x"1e",x"49"),
  1147 => (x"87",x"f5",x"da",x"c1"),
  1148 => (x"48",x"e0",x"f1",x"c2"),
  1149 => (x"49",x"c1",x"78",x"de"),
  1150 => (x"26",x"87",x"ca",x"d6"),
  1151 => (x"1e",x"87",x"fe",x"f6"),
  1152 => (x"cb",x"49",x"4a",x"71"),
  1153 => (x"d0",x"e2",x"c1",x"91"),
  1154 => (x"11",x"81",x"c8",x"81"),
  1155 => (x"e4",x"f1",x"c2",x"48"),
  1156 => (x"e4",x"f1",x"c2",x"58"),
  1157 => (x"c1",x"78",x"c0",x"48"),
  1158 => (x"87",x"e9",x"d5",x"49"),
  1159 => (x"c0",x"1e",x"4f",x"26"),
  1160 => (x"ca",x"c7",x"c1",x"49"),
  1161 => (x"1e",x"4f",x"26",x"87"),
  1162 => (x"d2",x"02",x"99",x"71"),
  1163 => (x"e5",x"e3",x"c1",x"87"),
  1164 => (x"f7",x"50",x"c0",x"48"),
  1165 => (x"ff",x"c7",x"c1",x"80"),
  1166 => (x"c9",x"e2",x"c1",x"40"),
  1167 => (x"c1",x"87",x"ce",x"78"),
  1168 => (x"c1",x"48",x"e1",x"e3"),
  1169 => (x"fc",x"78",x"c2",x"e2"),
  1170 => (x"de",x"c8",x"c1",x"80"),
  1171 => (x"0e",x"4f",x"26",x"78"),
  1172 => (x"0e",x"5c",x"5b",x"5e"),
  1173 => (x"cb",x"4a",x"4c",x"71"),
  1174 => (x"d0",x"e2",x"c1",x"92"),
  1175 => (x"49",x"a2",x"c8",x"82"),
  1176 => (x"97",x"4b",x"a2",x"c9"),
  1177 => (x"97",x"1e",x"4b",x"6b"),
  1178 => (x"ca",x"1e",x"49",x"69"),
  1179 => (x"c0",x"49",x"12",x"82"),
  1180 => (x"c0",x"87",x"eb",x"e7"),
  1181 => (x"87",x"cd",x"d4",x"49"),
  1182 => (x"c4",x"c1",x"49",x"74"),
  1183 => (x"8e",x"f8",x"87",x"cc"),
  1184 => (x"1e",x"87",x"f8",x"f4"),
  1185 => (x"4b",x"71",x"1e",x"73"),
  1186 => (x"87",x"c3",x"ff",x"49"),
  1187 => (x"fe",x"fe",x"49",x"73"),
  1188 => (x"87",x"e9",x"f4",x"87"),
  1189 => (x"71",x"1e",x"73",x"1e"),
  1190 => (x"4a",x"a3",x"c6",x"4b"),
  1191 => (x"c1",x"87",x"db",x"02"),
  1192 => (x"87",x"d6",x"02",x"8a"),
  1193 => (x"da",x"c1",x"02",x"8a"),
  1194 => (x"c0",x"02",x"8a",x"87"),
  1195 => (x"02",x"8a",x"87",x"fc"),
  1196 => (x"8a",x"87",x"e1",x"c0"),
  1197 => (x"c1",x"87",x"cb",x"02"),
  1198 => (x"49",x"c7",x"87",x"db"),
  1199 => (x"c1",x"87",x"c0",x"fd"),
  1200 => (x"f1",x"c2",x"87",x"de"),
  1201 => (x"c1",x"02",x"bf",x"e4"),
  1202 => (x"c1",x"48",x"87",x"cb"),
  1203 => (x"e8",x"f1",x"c2",x"88"),
  1204 => (x"87",x"c1",x"c1",x"58"),
  1205 => (x"bf",x"e8",x"f1",x"c2"),
  1206 => (x"87",x"f9",x"c0",x"02"),
  1207 => (x"bf",x"e4",x"f1",x"c2"),
  1208 => (x"c2",x"80",x"c1",x"48"),
  1209 => (x"c0",x"58",x"e8",x"f1"),
  1210 => (x"f1",x"c2",x"87",x"eb"),
  1211 => (x"c6",x"49",x"bf",x"e4"),
  1212 => (x"e8",x"f1",x"c2",x"89"),
  1213 => (x"a9",x"b7",x"c0",x"59"),
  1214 => (x"c2",x"87",x"da",x"03"),
  1215 => (x"c0",x"48",x"e4",x"f1"),
  1216 => (x"c2",x"87",x"d2",x"78"),
  1217 => (x"02",x"bf",x"e8",x"f1"),
  1218 => (x"f1",x"c2",x"87",x"cb"),
  1219 => (x"c6",x"48",x"bf",x"e4"),
  1220 => (x"e8",x"f1",x"c2",x"80"),
  1221 => (x"d1",x"49",x"c0",x"58"),
  1222 => (x"49",x"73",x"87",x"eb"),
  1223 => (x"87",x"ea",x"c1",x"c1"),
  1224 => (x"1e",x"87",x"da",x"f2"),
  1225 => (x"4b",x"71",x"1e",x"73"),
  1226 => (x"48",x"e0",x"f1",x"c2"),
  1227 => (x"49",x"c0",x"78",x"dd"),
  1228 => (x"73",x"87",x"d2",x"d1"),
  1229 => (x"d1",x"c1",x"c1",x"49"),
  1230 => (x"87",x"c1",x"f2",x"87"),
  1231 => (x"5c",x"5b",x"5e",x"0e"),
  1232 => (x"cc",x"4c",x"71",x"0e"),
  1233 => (x"4b",x"74",x"1e",x"66"),
  1234 => (x"e2",x"c1",x"93",x"cb"),
  1235 => (x"a3",x"c4",x"83",x"d0"),
  1236 => (x"fe",x"49",x"6a",x"4a"),
  1237 => (x"c1",x"87",x"e1",x"f5"),
  1238 => (x"c8",x"7b",x"fd",x"c6"),
  1239 => (x"66",x"d4",x"49",x"a3"),
  1240 => (x"49",x"a3",x"c9",x"51"),
  1241 => (x"ca",x"51",x"66",x"d8"),
  1242 => (x"66",x"dc",x"49",x"a3"),
  1243 => (x"ca",x"f1",x"26",x"51"),
  1244 => (x"5b",x"5e",x"0e",x"87"),
  1245 => (x"ff",x"0e",x"5d",x"5c"),
  1246 => (x"a6",x"dc",x"86",x"cc"),
  1247 => (x"48",x"a6",x"c8",x"59"),
  1248 => (x"80",x"c4",x"78",x"c0"),
  1249 => (x"78",x"66",x"c8",x"c1"),
  1250 => (x"78",x"c1",x"80",x"c4"),
  1251 => (x"78",x"c1",x"80",x"c4"),
  1252 => (x"48",x"e8",x"f1",x"c2"),
  1253 => (x"f1",x"c2",x"78",x"c1"),
  1254 => (x"de",x"48",x"bf",x"e0"),
  1255 => (x"87",x"cb",x"05",x"a8"),
  1256 => (x"70",x"87",x"cc",x"f3"),
  1257 => (x"59",x"a6",x"cc",x"49"),
  1258 => (x"e7",x"87",x"d6",x"ce"),
  1259 => (x"c4",x"e8",x"87",x"d2"),
  1260 => (x"87",x"ec",x"e6",x"87"),
  1261 => (x"fb",x"c0",x"4c",x"70"),
  1262 => (x"d8",x"c1",x"02",x"ac"),
  1263 => (x"05",x"66",x"d8",x"87"),
  1264 => (x"c0",x"87",x"ca",x"c1"),
  1265 => (x"1e",x"c1",x"1e",x"1e"),
  1266 => (x"1e",x"c3",x"e4",x"c1"),
  1267 => (x"eb",x"fd",x"49",x"c0"),
  1268 => (x"c0",x"86",x"d0",x"87"),
  1269 => (x"d9",x"02",x"ac",x"fb"),
  1270 => (x"66",x"c4",x"c1",x"87"),
  1271 => (x"6a",x"82",x"c4",x"4a"),
  1272 => (x"74",x"81",x"c7",x"49"),
  1273 => (x"d8",x"1e",x"c1",x"51"),
  1274 => (x"c8",x"49",x"6a",x"1e"),
  1275 => (x"87",x"d9",x"e7",x"81"),
  1276 => (x"c8",x"c1",x"86",x"c8"),
  1277 => (x"a8",x"c0",x"48",x"66"),
  1278 => (x"c8",x"87",x"c7",x"01"),
  1279 => (x"78",x"c1",x"48",x"a6"),
  1280 => (x"c8",x"c1",x"87",x"ce"),
  1281 => (x"88",x"c1",x"48",x"66"),
  1282 => (x"c3",x"58",x"a6",x"d0"),
  1283 => (x"87",x"e5",x"e6",x"87"),
  1284 => (x"c2",x"48",x"a6",x"d0"),
  1285 => (x"02",x"9c",x"74",x"78"),
  1286 => (x"c8",x"87",x"e2",x"cc"),
  1287 => (x"cc",x"c1",x"48",x"66"),
  1288 => (x"cc",x"03",x"a8",x"66"),
  1289 => (x"a6",x"dc",x"87",x"d7"),
  1290 => (x"e4",x"78",x"c0",x"48"),
  1291 => (x"4c",x"70",x"87",x"f2"),
  1292 => (x"dd",x"48",x"66",x"d8"),
  1293 => (x"87",x"c6",x"05",x"a8"),
  1294 => (x"d8",x"48",x"a6",x"dc"),
  1295 => (x"d0",x"c1",x"78",x"66"),
  1296 => (x"e8",x"c0",x"05",x"ac"),
  1297 => (x"87",x"d8",x"e4",x"87"),
  1298 => (x"70",x"87",x"d5",x"e4"),
  1299 => (x"ac",x"ec",x"c0",x"4c"),
  1300 => (x"e5",x"87",x"c5",x"05"),
  1301 => (x"4c",x"70",x"87",x"df"),
  1302 => (x"05",x"ac",x"d0",x"c1"),
  1303 => (x"66",x"d4",x"87",x"c8"),
  1304 => (x"d8",x"80",x"c1",x"48"),
  1305 => (x"d0",x"c1",x"58",x"a6"),
  1306 => (x"d8",x"ff",x"02",x"ac"),
  1307 => (x"a6",x"e0",x"c0",x"87"),
  1308 => (x"78",x"66",x"d8",x"48"),
  1309 => (x"c0",x"48",x"66",x"dc"),
  1310 => (x"05",x"a8",x"66",x"e0"),
  1311 => (x"c4",x"87",x"d0",x"ca"),
  1312 => (x"f0",x"c0",x"48",x"a6"),
  1313 => (x"80",x"e0",x"c0",x"78"),
  1314 => (x"c4",x"78",x"66",x"d0"),
  1315 => (x"c4",x"78",x"c0",x"80"),
  1316 => (x"74",x"78",x"c0",x"80"),
  1317 => (x"8d",x"fb",x"c0",x"4d"),
  1318 => (x"87",x"cc",x"c9",x"02"),
  1319 => (x"db",x"02",x"8d",x"c9"),
  1320 => (x"02",x"8d",x"c2",x"87"),
  1321 => (x"c9",x"87",x"cd",x"c1"),
  1322 => (x"d1",x"c4",x"02",x"8d"),
  1323 => (x"02",x"8d",x"c4",x"87"),
  1324 => (x"c1",x"87",x"ce",x"c1"),
  1325 => (x"c5",x"c4",x"02",x"8d"),
  1326 => (x"87",x"e6",x"c8",x"87"),
  1327 => (x"cb",x"49",x"66",x"c8"),
  1328 => (x"66",x"c4",x"c1",x"91"),
  1329 => (x"4a",x"a1",x"c4",x"81"),
  1330 => (x"1e",x"71",x"7e",x"6a"),
  1331 => (x"48",x"f8",x"dd",x"c1"),
  1332 => (x"cc",x"49",x"66",x"c4"),
  1333 => (x"41",x"20",x"4a",x"a1"),
  1334 => (x"ff",x"05",x"aa",x"71"),
  1335 => (x"51",x"10",x"87",x"f8"),
  1336 => (x"cc",x"c1",x"49",x"26"),
  1337 => (x"cc",x"e3",x"79",x"e3"),
  1338 => (x"c0",x"4c",x"70",x"87"),
  1339 => (x"c1",x"48",x"a6",x"ec"),
  1340 => (x"87",x"f4",x"c7",x"78"),
  1341 => (x"c0",x"48",x"a6",x"c4"),
  1342 => (x"48",x"66",x"d0",x"78"),
  1343 => (x"a6",x"d4",x"80",x"c1"),
  1344 => (x"87",x"dc",x"e1",x"58"),
  1345 => (x"ec",x"c0",x"4c",x"70"),
  1346 => (x"87",x"d4",x"02",x"ac"),
  1347 => (x"c0",x"02",x"66",x"c4"),
  1348 => (x"a6",x"c8",x"87",x"c5"),
  1349 => (x"74",x"87",x"c9",x"5c"),
  1350 => (x"88",x"f0",x"c0",x"48"),
  1351 => (x"58",x"a6",x"e8",x"c0"),
  1352 => (x"02",x"ac",x"ec",x"c0"),
  1353 => (x"f7",x"e0",x"87",x"cc"),
  1354 => (x"c0",x"4c",x"70",x"87"),
  1355 => (x"ff",x"05",x"ac",x"ec"),
  1356 => (x"66",x"c4",x"87",x"f4"),
  1357 => (x"49",x"66",x"d8",x"1e"),
  1358 => (x"66",x"ec",x"c0",x"1e"),
  1359 => (x"c3",x"e4",x"c1",x"1e"),
  1360 => (x"49",x"66",x"d8",x"1e"),
  1361 => (x"c0",x"87",x"f5",x"f7"),
  1362 => (x"c0",x"1e",x"ca",x"1e"),
  1363 => (x"cb",x"49",x"66",x"e0"),
  1364 => (x"66",x"dc",x"c1",x"91"),
  1365 => (x"48",x"a6",x"d8",x"81"),
  1366 => (x"d8",x"78",x"a1",x"c4"),
  1367 => (x"e1",x"49",x"bf",x"66"),
  1368 => (x"86",x"d8",x"87",x"e7"),
  1369 => (x"06",x"a8",x"b7",x"c0"),
  1370 => (x"c1",x"87",x"ca",x"c1"),
  1371 => (x"c8",x"1e",x"de",x"1e"),
  1372 => (x"e1",x"49",x"bf",x"66"),
  1373 => (x"86",x"c8",x"87",x"d3"),
  1374 => (x"c0",x"48",x"49",x"70"),
  1375 => (x"e8",x"c0",x"88",x"08"),
  1376 => (x"b7",x"c0",x"58",x"a6"),
  1377 => (x"ec",x"c0",x"06",x"a8"),
  1378 => (x"66",x"e4",x"c0",x"87"),
  1379 => (x"a8",x"b7",x"dd",x"48"),
  1380 => (x"87",x"e1",x"c0",x"03"),
  1381 => (x"c0",x"49",x"bf",x"6e"),
  1382 => (x"c0",x"81",x"66",x"e4"),
  1383 => (x"e4",x"c0",x"51",x"e0"),
  1384 => (x"81",x"c1",x"49",x"66"),
  1385 => (x"c2",x"81",x"bf",x"6e"),
  1386 => (x"e4",x"c0",x"51",x"c1"),
  1387 => (x"81",x"c2",x"49",x"66"),
  1388 => (x"c0",x"81",x"bf",x"6e"),
  1389 => (x"a6",x"ec",x"c0",x"51"),
  1390 => (x"c4",x"78",x"c1",x"48"),
  1391 => (x"f7",x"e1",x"87",x"ea"),
  1392 => (x"a6",x"e8",x"c0",x"87"),
  1393 => (x"87",x"f0",x"e1",x"58"),
  1394 => (x"58",x"a6",x"f0",x"c0"),
  1395 => (x"05",x"a8",x"ec",x"c0"),
  1396 => (x"a6",x"87",x"c9",x"c0"),
  1397 => (x"66",x"e4",x"c0",x"48"),
  1398 => (x"87",x"c4",x"c0",x"78"),
  1399 => (x"87",x"c0",x"de",x"ff"),
  1400 => (x"cb",x"49",x"66",x"c8"),
  1401 => (x"66",x"c4",x"c1",x"91"),
  1402 => (x"c8",x"80",x"71",x"48"),
  1403 => (x"66",x"c4",x"58",x"a6"),
  1404 => (x"c4",x"82",x"c8",x"4a"),
  1405 => (x"81",x"ca",x"49",x"66"),
  1406 => (x"51",x"66",x"e4",x"c0"),
  1407 => (x"49",x"66",x"ec",x"c0"),
  1408 => (x"e4",x"c0",x"81",x"c1"),
  1409 => (x"48",x"c1",x"89",x"66"),
  1410 => (x"49",x"70",x"30",x"71"),
  1411 => (x"97",x"71",x"89",x"c1"),
  1412 => (x"d5",x"f5",x"c2",x"7a"),
  1413 => (x"e4",x"c0",x"49",x"bf"),
  1414 => (x"6a",x"97",x"29",x"66"),
  1415 => (x"98",x"71",x"48",x"4a"),
  1416 => (x"58",x"a6",x"f4",x"c0"),
  1417 => (x"c4",x"49",x"66",x"c4"),
  1418 => (x"c0",x"7e",x"69",x"81"),
  1419 => (x"dc",x"48",x"66",x"e0"),
  1420 => (x"c0",x"02",x"a8",x"66"),
  1421 => (x"a6",x"dc",x"87",x"c8"),
  1422 => (x"c0",x"78",x"c0",x"48"),
  1423 => (x"a6",x"dc",x"87",x"c5"),
  1424 => (x"dc",x"78",x"c1",x"48"),
  1425 => (x"e0",x"c0",x"1e",x"66"),
  1426 => (x"49",x"66",x"c8",x"1e"),
  1427 => (x"87",x"f9",x"dd",x"ff"),
  1428 => (x"4c",x"70",x"86",x"c8"),
  1429 => (x"06",x"ac",x"b7",x"c0"),
  1430 => (x"6e",x"87",x"d6",x"c1"),
  1431 => (x"70",x"80",x"74",x"48"),
  1432 => (x"49",x"e0",x"c0",x"7e"),
  1433 => (x"4b",x"6e",x"89",x"74"),
  1434 => (x"4a",x"f5",x"dd",x"c1"),
  1435 => (x"f7",x"e8",x"fe",x"71"),
  1436 => (x"c2",x"48",x"6e",x"87"),
  1437 => (x"c0",x"7e",x"70",x"80"),
  1438 => (x"c1",x"48",x"66",x"e8"),
  1439 => (x"a6",x"ec",x"c0",x"80"),
  1440 => (x"66",x"f0",x"c0",x"58"),
  1441 => (x"70",x"81",x"c1",x"49"),
  1442 => (x"c5",x"c0",x"02",x"a9"),
  1443 => (x"c0",x"4d",x"c0",x"87"),
  1444 => (x"4d",x"c1",x"87",x"c2"),
  1445 => (x"a4",x"c2",x"1e",x"75"),
  1446 => (x"48",x"e0",x"c0",x"49"),
  1447 => (x"49",x"70",x"88",x"71"),
  1448 => (x"49",x"66",x"c8",x"1e"),
  1449 => (x"87",x"e1",x"dc",x"ff"),
  1450 => (x"b7",x"c0",x"86",x"c8"),
  1451 => (x"c6",x"ff",x"01",x"a8"),
  1452 => (x"66",x"e8",x"c0",x"87"),
  1453 => (x"87",x"d3",x"c0",x"02"),
  1454 => (x"c9",x"49",x"66",x"c4"),
  1455 => (x"66",x"e8",x"c0",x"81"),
  1456 => (x"48",x"66",x"c4",x"51"),
  1457 => (x"78",x"cf",x"c9",x"c1"),
  1458 => (x"c4",x"87",x"ce",x"c0"),
  1459 => (x"81",x"c9",x"49",x"66"),
  1460 => (x"66",x"c4",x"51",x"c2"),
  1461 => (x"c3",x"ca",x"c1",x"48"),
  1462 => (x"a6",x"ec",x"c0",x"78"),
  1463 => (x"c0",x"78",x"c1",x"48"),
  1464 => (x"db",x"ff",x"87",x"c6"),
  1465 => (x"4c",x"70",x"87",x"cf"),
  1466 => (x"02",x"66",x"ec",x"c0"),
  1467 => (x"c8",x"87",x"f5",x"c0"),
  1468 => (x"66",x"cc",x"48",x"66"),
  1469 => (x"cb",x"c0",x"04",x"a8"),
  1470 => (x"48",x"66",x"c8",x"87"),
  1471 => (x"a6",x"cc",x"80",x"c1"),
  1472 => (x"87",x"e0",x"c0",x"58"),
  1473 => (x"c1",x"48",x"66",x"cc"),
  1474 => (x"58",x"a6",x"d0",x"88"),
  1475 => (x"c1",x"87",x"d5",x"c0"),
  1476 => (x"c0",x"05",x"ac",x"c6"),
  1477 => (x"66",x"d0",x"87",x"c8"),
  1478 => (x"d4",x"80",x"c1",x"48"),
  1479 => (x"da",x"ff",x"58",x"a6"),
  1480 => (x"4c",x"70",x"87",x"d3"),
  1481 => (x"c1",x"48",x"66",x"d4"),
  1482 => (x"58",x"a6",x"d8",x"80"),
  1483 => (x"c0",x"02",x"9c",x"74"),
  1484 => (x"66",x"c8",x"87",x"cb"),
  1485 => (x"66",x"cc",x"c1",x"48"),
  1486 => (x"e9",x"f3",x"04",x"a8"),
  1487 => (x"eb",x"d9",x"ff",x"87"),
  1488 => (x"48",x"66",x"c8",x"87"),
  1489 => (x"c0",x"03",x"a8",x"c7"),
  1490 => (x"f1",x"c2",x"87",x"e5"),
  1491 => (x"78",x"c0",x"48",x"e8"),
  1492 => (x"cb",x"49",x"66",x"c8"),
  1493 => (x"66",x"c4",x"c1",x"91"),
  1494 => (x"4a",x"a1",x"c4",x"81"),
  1495 => (x"52",x"c0",x"4a",x"6a"),
  1496 => (x"48",x"66",x"c8",x"79"),
  1497 => (x"a6",x"cc",x"80",x"c1"),
  1498 => (x"04",x"a8",x"c7",x"58"),
  1499 => (x"ff",x"87",x"db",x"ff"),
  1500 => (x"c4",x"e1",x"8e",x"cc"),
  1501 => (x"00",x"20",x"3a",x"87"),
  1502 => (x"20",x"50",x"49",x"44"),
  1503 => (x"74",x"69",x"77",x"53"),
  1504 => (x"73",x"65",x"68",x"63"),
  1505 => (x"1e",x"73",x"1e",x"00"),
  1506 => (x"02",x"9b",x"4b",x"71"),
  1507 => (x"f1",x"c2",x"87",x"c6"),
  1508 => (x"78",x"c0",x"48",x"e4"),
  1509 => (x"f1",x"c2",x"1e",x"c7"),
  1510 => (x"1e",x"49",x"bf",x"e4"),
  1511 => (x"1e",x"d0",x"e2",x"c1"),
  1512 => (x"bf",x"e0",x"f1",x"c2"),
  1513 => (x"87",x"c9",x"ef",x"49"),
  1514 => (x"f1",x"c2",x"86",x"cc"),
  1515 => (x"e9",x"49",x"bf",x"e0"),
  1516 => (x"9b",x"73",x"87",x"f5"),
  1517 => (x"c1",x"87",x"c8",x"02"),
  1518 => (x"c0",x"49",x"d0",x"e2"),
  1519 => (x"ff",x"87",x"dd",x"f0"),
  1520 => (x"1e",x"87",x"fa",x"df"),
  1521 => (x"4b",x"c0",x"1e",x"73"),
  1522 => (x"48",x"f4",x"e2",x"c2"),
  1523 => (x"e3",x"c1",x"50",x"c0"),
  1524 => (x"c0",x"49",x"bf",x"f3"),
  1525 => (x"70",x"87",x"e5",x"fe"),
  1526 => (x"87",x"c4",x"05",x"98"),
  1527 => (x"4b",x"e6",x"df",x"c1"),
  1528 => (x"df",x"ff",x"48",x"73"),
  1529 => (x"4f",x"52",x"87",x"d7"),
  1530 => (x"6f",x"6c",x"20",x"4d"),
  1531 => (x"6e",x"69",x"64",x"61"),
  1532 => (x"61",x"66",x"20",x"67"),
  1533 => (x"64",x"65",x"6c",x"69"),
  1534 => (x"e5",x"c7",x"1e",x"00"),
  1535 => (x"fe",x"49",x"c1",x"87"),
  1536 => (x"ea",x"fe",x"87",x"c3"),
  1537 => (x"98",x"70",x"87",x"ec"),
  1538 => (x"fe",x"87",x"cd",x"02"),
  1539 => (x"70",x"87",x"c7",x"f2"),
  1540 => (x"87",x"c4",x"02",x"98"),
  1541 => (x"87",x"c2",x"4a",x"c1"),
  1542 => (x"9a",x"72",x"4a",x"c0"),
  1543 => (x"c0",x"87",x"ce",x"05"),
  1544 => (x"cd",x"e1",x"c1",x"1e"),
  1545 => (x"d1",x"fb",x"c0",x"49"),
  1546 => (x"fe",x"86",x"c4",x"87"),
  1547 => (x"ed",x"c2",x"c1",x"87"),
  1548 => (x"c1",x"1e",x"c0",x"87"),
  1549 => (x"c0",x"49",x"d8",x"e1"),
  1550 => (x"c0",x"87",x"ff",x"fa"),
  1551 => (x"87",x"c3",x"fe",x"1e"),
  1552 => (x"fa",x"c0",x"49",x"70"),
  1553 => (x"d8",x"c3",x"87",x"f4"),
  1554 => (x"26",x"8e",x"f8",x"87"),
  1555 => (x"20",x"44",x"53",x"4f"),
  1556 => (x"6c",x"69",x"61",x"66"),
  1557 => (x"00",x"2e",x"64",x"65"),
  1558 => (x"74",x"6f",x"6f",x"42"),
  1559 => (x"2e",x"67",x"6e",x"69"),
  1560 => (x"1e",x"00",x"2e",x"2e"),
  1561 => (x"87",x"d5",x"f2",x"c0"),
  1562 => (x"4f",x"26",x"87",x"fa"),
  1563 => (x"e4",x"f1",x"c2",x"1e"),
  1564 => (x"c2",x"78",x"c0",x"48"),
  1565 => (x"c0",x"48",x"e0",x"f1"),
  1566 => (x"87",x"fd",x"fd",x"78"),
  1567 => (x"48",x"c0",x"87",x"e5"),
  1568 => (x"20",x"80",x"4f",x"26"),
  1569 => (x"74",x"69",x"78",x"45"),
  1570 => (x"42",x"20",x"80",x"00"),
  1571 => (x"00",x"6b",x"63",x"61"),
  1572 => (x"00",x"00",x"11",x"ff"),
  1573 => (x"00",x"00",x"2c",x"79"),
  1574 => (x"ff",x"00",x"00",x"00"),
  1575 => (x"97",x"00",x"00",x"11"),
  1576 => (x"00",x"00",x"00",x"2c"),
  1577 => (x"11",x"ff",x"00",x"00"),
  1578 => (x"2c",x"b5",x"00",x"00"),
  1579 => (x"00",x"00",x"00",x"00"),
  1580 => (x"00",x"11",x"ff",x"00"),
  1581 => (x"00",x"2c",x"d3",x"00"),
  1582 => (x"00",x"00",x"00",x"00"),
  1583 => (x"00",x"00",x"11",x"ff"),
  1584 => (x"00",x"00",x"2c",x"f1"),
  1585 => (x"ff",x"00",x"00",x"00"),
  1586 => (x"0f",x"00",x"00",x"11"),
  1587 => (x"00",x"00",x"00",x"2d"),
  1588 => (x"11",x"ff",x"00",x"00"),
  1589 => (x"2d",x"2d",x"00",x"00"),
  1590 => (x"00",x"00",x"00",x"00"),
  1591 => (x"00",x"11",x"ff",x"00"),
  1592 => (x"00",x"00",x"00",x"00"),
  1593 => (x"00",x"00",x"00",x"00"),
  1594 => (x"00",x"00",x"12",x"94"),
  1595 => (x"00",x"00",x"00",x"00"),
  1596 => (x"f7",x"00",x"00",x"00"),
  1597 => (x"4d",x"00",x"00",x"18"),
  1598 => (x"20",x"55",x"4e",x"45"),
  1599 => (x"52",x"20",x"20",x"20"),
  1600 => (x"4c",x"00",x"4d",x"4f"),
  1601 => (x"20",x"64",x"61",x"6f"),
  1602 => (x"1e",x"00",x"2e",x"2a"),
  1603 => (x"c0",x"48",x"f0",x"fe"),
  1604 => (x"79",x"09",x"cd",x"78"),
  1605 => (x"1e",x"4f",x"26",x"09"),
  1606 => (x"bf",x"f0",x"fe",x"1e"),
  1607 => (x"26",x"26",x"48",x"7e"),
  1608 => (x"f0",x"fe",x"1e",x"4f"),
  1609 => (x"26",x"78",x"c1",x"48"),
  1610 => (x"f0",x"fe",x"1e",x"4f"),
  1611 => (x"26",x"78",x"c0",x"48"),
  1612 => (x"4a",x"71",x"1e",x"4f"),
  1613 => (x"26",x"52",x"52",x"c0"),
  1614 => (x"5b",x"5e",x"0e",x"4f"),
  1615 => (x"f4",x"0e",x"5d",x"5c"),
  1616 => (x"97",x"4d",x"71",x"86"),
  1617 => (x"a5",x"c1",x"7e",x"6d"),
  1618 => (x"48",x"6c",x"97",x"4c"),
  1619 => (x"6e",x"58",x"a6",x"c8"),
  1620 => (x"a8",x"66",x"c4",x"48"),
  1621 => (x"ff",x"87",x"c5",x"05"),
  1622 => (x"87",x"e6",x"c0",x"48"),
  1623 => (x"c2",x"87",x"ca",x"ff"),
  1624 => (x"6c",x"97",x"49",x"a5"),
  1625 => (x"4b",x"a3",x"71",x"4b"),
  1626 => (x"97",x"4b",x"6b",x"97"),
  1627 => (x"48",x"6e",x"7e",x"6c"),
  1628 => (x"a6",x"c8",x"80",x"c1"),
  1629 => (x"cc",x"98",x"c7",x"58"),
  1630 => (x"97",x"70",x"58",x"a6"),
  1631 => (x"87",x"e1",x"fe",x"7c"),
  1632 => (x"8e",x"f4",x"48",x"73"),
  1633 => (x"4c",x"26",x"4d",x"26"),
  1634 => (x"4f",x"26",x"4b",x"26"),
  1635 => (x"5c",x"5b",x"5e",x"0e"),
  1636 => (x"71",x"86",x"f4",x"0e"),
  1637 => (x"4a",x"66",x"d8",x"4c"),
  1638 => (x"c2",x"9a",x"ff",x"c3"),
  1639 => (x"6c",x"97",x"4b",x"a4"),
  1640 => (x"49",x"a1",x"73",x"49"),
  1641 => (x"6c",x"97",x"51",x"72"),
  1642 => (x"c1",x"48",x"6e",x"7e"),
  1643 => (x"58",x"a6",x"c8",x"80"),
  1644 => (x"a6",x"cc",x"98",x"c7"),
  1645 => (x"f4",x"54",x"70",x"58"),
  1646 => (x"87",x"ca",x"ff",x"8e"),
  1647 => (x"e8",x"fd",x"1e",x"1e"),
  1648 => (x"4a",x"bf",x"e0",x"87"),
  1649 => (x"c0",x"e0",x"c0",x"49"),
  1650 => (x"87",x"cb",x"02",x"99"),
  1651 => (x"f5",x"c2",x"1e",x"72"),
  1652 => (x"f7",x"fe",x"49",x"cb"),
  1653 => (x"fc",x"86",x"c4",x"87"),
  1654 => (x"7e",x"70",x"87",x"fd"),
  1655 => (x"26",x"87",x"c2",x"fd"),
  1656 => (x"c2",x"1e",x"4f",x"26"),
  1657 => (x"fd",x"49",x"cb",x"f5"),
  1658 => (x"e6",x"c1",x"87",x"c7"),
  1659 => (x"da",x"fc",x"49",x"fc"),
  1660 => (x"87",x"d9",x"c5",x"87"),
  1661 => (x"5e",x"0e",x"4f",x"26"),
  1662 => (x"0e",x"5d",x"5c",x"5b"),
  1663 => (x"bf",x"de",x"f6",x"c2"),
  1664 => (x"ca",x"e9",x"c1",x"4a"),
  1665 => (x"72",x"4c",x"49",x"bf"),
  1666 => (x"fc",x"4d",x"71",x"bc"),
  1667 => (x"4b",x"c0",x"87",x"db"),
  1668 => (x"99",x"d0",x"49",x"74"),
  1669 => (x"75",x"87",x"d5",x"02"),
  1670 => (x"71",x"99",x"d0",x"49"),
  1671 => (x"c1",x"1e",x"c0",x"1e"),
  1672 => (x"73",x"4a",x"dc",x"ef"),
  1673 => (x"c0",x"49",x"12",x"82"),
  1674 => (x"86",x"c8",x"87",x"e4"),
  1675 => (x"83",x"2d",x"2c",x"c1"),
  1676 => (x"ff",x"04",x"ab",x"c8"),
  1677 => (x"e8",x"fb",x"87",x"da"),
  1678 => (x"ca",x"e9",x"c1",x"87"),
  1679 => (x"de",x"f6",x"c2",x"48"),
  1680 => (x"4d",x"26",x"78",x"bf"),
  1681 => (x"4b",x"26",x"4c",x"26"),
  1682 => (x"00",x"00",x"4f",x"26"),
  1683 => (x"ff",x"1e",x"00",x"00"),
  1684 => (x"e1",x"c8",x"48",x"d0"),
  1685 => (x"48",x"d4",x"ff",x"78"),
  1686 => (x"66",x"c4",x"78",x"c5"),
  1687 => (x"c3",x"87",x"c3",x"02"),
  1688 => (x"66",x"c8",x"78",x"e0"),
  1689 => (x"ff",x"87",x"c6",x"02"),
  1690 => (x"f0",x"c3",x"48",x"d4"),
  1691 => (x"48",x"d4",x"ff",x"78"),
  1692 => (x"d0",x"ff",x"78",x"71"),
  1693 => (x"78",x"e1",x"c8",x"48"),
  1694 => (x"26",x"78",x"e0",x"c0"),
  1695 => (x"5b",x"5e",x"0e",x"4f"),
  1696 => (x"4c",x"71",x"0e",x"5c"),
  1697 => (x"49",x"cb",x"f5",x"c2"),
  1698 => (x"70",x"87",x"ee",x"fa"),
  1699 => (x"aa",x"b7",x"c0",x"4a"),
  1700 => (x"87",x"e3",x"c2",x"04"),
  1701 => (x"05",x"aa",x"e0",x"c3"),
  1702 => (x"ed",x"c1",x"87",x"c9"),
  1703 => (x"78",x"c1",x"48",x"c0"),
  1704 => (x"c3",x"87",x"d4",x"c2"),
  1705 => (x"c9",x"05",x"aa",x"f0"),
  1706 => (x"fc",x"ec",x"c1",x"87"),
  1707 => (x"c1",x"78",x"c1",x"48"),
  1708 => (x"ed",x"c1",x"87",x"f5"),
  1709 => (x"c7",x"02",x"bf",x"c0"),
  1710 => (x"c2",x"4b",x"72",x"87"),
  1711 => (x"87",x"c2",x"b3",x"c0"),
  1712 => (x"9c",x"74",x"4b",x"72"),
  1713 => (x"c1",x"87",x"d1",x"05"),
  1714 => (x"1e",x"bf",x"fc",x"ec"),
  1715 => (x"bf",x"c0",x"ed",x"c1"),
  1716 => (x"fd",x"49",x"72",x"1e"),
  1717 => (x"86",x"c8",x"87",x"f8"),
  1718 => (x"bf",x"fc",x"ec",x"c1"),
  1719 => (x"87",x"e0",x"c0",x"02"),
  1720 => (x"b7",x"c4",x"49",x"73"),
  1721 => (x"ee",x"c1",x"91",x"29"),
  1722 => (x"4a",x"73",x"81",x"dc"),
  1723 => (x"92",x"c2",x"9a",x"cf"),
  1724 => (x"30",x"72",x"48",x"c1"),
  1725 => (x"ba",x"ff",x"4a",x"70"),
  1726 => (x"98",x"69",x"48",x"72"),
  1727 => (x"87",x"db",x"79",x"70"),
  1728 => (x"b7",x"c4",x"49",x"73"),
  1729 => (x"ee",x"c1",x"91",x"29"),
  1730 => (x"4a",x"73",x"81",x"dc"),
  1731 => (x"92",x"c2",x"9a",x"cf"),
  1732 => (x"30",x"72",x"48",x"c3"),
  1733 => (x"69",x"48",x"4a",x"70"),
  1734 => (x"c1",x"79",x"70",x"b0"),
  1735 => (x"c0",x"48",x"c0",x"ed"),
  1736 => (x"fc",x"ec",x"c1",x"78"),
  1737 => (x"c2",x"78",x"c0",x"48"),
  1738 => (x"f8",x"49",x"cb",x"f5"),
  1739 => (x"4a",x"70",x"87",x"cb"),
  1740 => (x"03",x"aa",x"b7",x"c0"),
  1741 => (x"c0",x"87",x"dd",x"fd"),
  1742 => (x"87",x"c8",x"fc",x"48"),
  1743 => (x"00",x"00",x"00",x"00"),
  1744 => (x"00",x"00",x"00",x"00"),
  1745 => (x"49",x"4a",x"71",x"1e"),
  1746 => (x"26",x"87",x"f2",x"fc"),
  1747 => (x"4a",x"c0",x"1e",x"4f"),
  1748 => (x"91",x"c4",x"49",x"72"),
  1749 => (x"81",x"dc",x"ee",x"c1"),
  1750 => (x"82",x"c1",x"79",x"c0"),
  1751 => (x"04",x"aa",x"b7",x"d0"),
  1752 => (x"4f",x"26",x"87",x"ee"),
  1753 => (x"5c",x"5b",x"5e",x"0e"),
  1754 => (x"4d",x"71",x"0e",x"5d"),
  1755 => (x"75",x"87",x"fa",x"f6"),
  1756 => (x"2a",x"b7",x"c4",x"4a"),
  1757 => (x"dc",x"ee",x"c1",x"92"),
  1758 => (x"cf",x"4c",x"75",x"82"),
  1759 => (x"6a",x"94",x"c2",x"9c"),
  1760 => (x"2b",x"74",x"4b",x"49"),
  1761 => (x"48",x"c2",x"9b",x"c3"),
  1762 => (x"4c",x"70",x"30",x"74"),
  1763 => (x"48",x"74",x"bc",x"ff"),
  1764 => (x"7a",x"70",x"98",x"71"),
  1765 => (x"73",x"87",x"ca",x"f6"),
  1766 => (x"87",x"e6",x"fa",x"48"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"25",x"26",x"1e",x"16"),
  1784 => (x"3e",x"3d",x"36",x"2e"),
  1785 => (x"48",x"d0",x"ff",x"1e"),
  1786 => (x"71",x"78",x"e1",x"c8"),
  1787 => (x"08",x"d4",x"ff",x"48"),
  1788 => (x"48",x"66",x"c4",x"78"),
  1789 => (x"78",x"08",x"d4",x"ff"),
  1790 => (x"71",x"1e",x"4f",x"26"),
  1791 => (x"49",x"66",x"c4",x"4a"),
  1792 => (x"ff",x"49",x"72",x"1e"),
  1793 => (x"d0",x"ff",x"87",x"de"),
  1794 => (x"78",x"e0",x"c0",x"48"),
  1795 => (x"1e",x"4f",x"26",x"26"),
  1796 => (x"66",x"c4",x"4a",x"71"),
  1797 => (x"a2",x"e0",x"c1",x"1e"),
  1798 => (x"87",x"c8",x"ff",x"49"),
  1799 => (x"c8",x"49",x"66",x"c8"),
  1800 => (x"d4",x"ff",x"29",x"b7"),
  1801 => (x"ff",x"78",x"71",x"48"),
  1802 => (x"e0",x"c0",x"48",x"d0"),
  1803 => (x"4f",x"26",x"26",x"78"),
  1804 => (x"4a",x"d4",x"ff",x"1e"),
  1805 => (x"ff",x"7a",x"ff",x"c3"),
  1806 => (x"e1",x"c8",x"48",x"d0"),
  1807 => (x"c2",x"7a",x"de",x"78"),
  1808 => (x"7a",x"bf",x"d5",x"f5"),
  1809 => (x"28",x"c8",x"48",x"49"),
  1810 => (x"48",x"71",x"7a",x"70"),
  1811 => (x"7a",x"70",x"28",x"d0"),
  1812 => (x"28",x"d8",x"48",x"71"),
  1813 => (x"d0",x"ff",x"7a",x"70"),
  1814 => (x"78",x"e0",x"c0",x"48"),
  1815 => (x"5e",x"0e",x"4f",x"26"),
  1816 => (x"0e",x"5d",x"5c",x"5b"),
  1817 => (x"f5",x"c2",x"4c",x"71"),
  1818 => (x"4b",x"4d",x"bf",x"d5"),
  1819 => (x"66",x"d0",x"2b",x"74"),
  1820 => (x"d4",x"83",x"c1",x"9b"),
  1821 => (x"c2",x"04",x"ab",x"66"),
  1822 => (x"74",x"4b",x"c0",x"87"),
  1823 => (x"49",x"66",x"d0",x"4a"),
  1824 => (x"b9",x"ff",x"31",x"72"),
  1825 => (x"48",x"73",x"99",x"75"),
  1826 => (x"4a",x"70",x"30",x"72"),
  1827 => (x"c2",x"b0",x"71",x"48"),
  1828 => (x"fe",x"58",x"d9",x"f5"),
  1829 => (x"4d",x"26",x"87",x"da"),
  1830 => (x"4b",x"26",x"4c",x"26"),
  1831 => (x"5e",x"0e",x"4f",x"26"),
  1832 => (x"0e",x"5d",x"5c",x"5b"),
  1833 => (x"c2",x"4c",x"71",x"1e"),
  1834 => (x"c0",x"4b",x"d9",x"f5"),
  1835 => (x"49",x"f4",x"c0",x"4a"),
  1836 => (x"87",x"d1",x"d0",x"fe"),
  1837 => (x"f5",x"c2",x"1e",x"74"),
  1838 => (x"ec",x"fe",x"49",x"d9"),
  1839 => (x"86",x"c4",x"87",x"e4"),
  1840 => (x"c0",x"02",x"98",x"70"),
  1841 => (x"1e",x"c4",x"87",x"ea"),
  1842 => (x"c2",x"1e",x"4d",x"a6"),
  1843 => (x"fe",x"49",x"d9",x"f5"),
  1844 => (x"c8",x"87",x"d5",x"f2"),
  1845 => (x"02",x"98",x"70",x"86"),
  1846 => (x"4a",x"75",x"87",x"d6"),
  1847 => (x"49",x"e6",x"f4",x"c1"),
  1848 => (x"ce",x"fe",x"4b",x"c4"),
  1849 => (x"98",x"70",x"87",x"c4"),
  1850 => (x"c0",x"87",x"ca",x"02"),
  1851 => (x"87",x"ed",x"c0",x"48"),
  1852 => (x"e8",x"c0",x"48",x"c0"),
  1853 => (x"87",x"f3",x"c0",x"87"),
  1854 => (x"70",x"87",x"c4",x"c1"),
  1855 => (x"87",x"c8",x"02",x"98"),
  1856 => (x"70",x"87",x"fc",x"c0"),
  1857 => (x"87",x"f8",x"05",x"98"),
  1858 => (x"bf",x"f9",x"f5",x"c2"),
  1859 => (x"c2",x"87",x"cc",x"02"),
  1860 => (x"c2",x"48",x"d5",x"f5"),
  1861 => (x"78",x"bf",x"f9",x"f5"),
  1862 => (x"c1",x"87",x"d5",x"fc"),
  1863 => (x"4d",x"26",x"26",x"48"),
  1864 => (x"4b",x"26",x"4c",x"26"),
  1865 => (x"41",x"5b",x"4f",x"26"),
  1866 => (x"1e",x"00",x"43",x"52"),
  1867 => (x"f5",x"c2",x"1e",x"c0"),
  1868 => (x"ef",x"fe",x"49",x"d9"),
  1869 => (x"f5",x"c2",x"87",x"cb"),
  1870 => (x"78",x"c0",x"48",x"f1"),
  1871 => (x"0e",x"4f",x"26",x"26"),
  1872 => (x"5d",x"5c",x"5b",x"5e"),
  1873 => (x"c4",x"86",x"f4",x"0e"),
  1874 => (x"78",x"c0",x"48",x"a6"),
  1875 => (x"bf",x"f1",x"f5",x"c2"),
  1876 => (x"a8",x"b7",x"c3",x"48"),
  1877 => (x"c2",x"87",x"d1",x"03"),
  1878 => (x"48",x"bf",x"f1",x"f5"),
  1879 => (x"f5",x"c2",x"80",x"c1"),
  1880 => (x"fb",x"c0",x"58",x"f5"),
  1881 => (x"87",x"e2",x"c6",x"48"),
  1882 => (x"49",x"d9",x"f5",x"c2"),
  1883 => (x"87",x"cc",x"f4",x"fe"),
  1884 => (x"f5",x"c2",x"4c",x"70"),
  1885 => (x"c3",x"4a",x"bf",x"f1"),
  1886 => (x"87",x"d8",x"02",x"8a"),
  1887 => (x"c5",x"02",x"8a",x"c1"),
  1888 => (x"02",x"8a",x"87",x"cb"),
  1889 => (x"8a",x"87",x"f6",x"c2"),
  1890 => (x"87",x"cd",x"c1",x"02"),
  1891 => (x"e2",x"c3",x"02",x"8a"),
  1892 => (x"87",x"e1",x"c5",x"87"),
  1893 => (x"4a",x"75",x"4d",x"c0"),
  1894 => (x"fc",x"c1",x"92",x"c4"),
  1895 => (x"f5",x"c2",x"82",x"e8"),
  1896 => (x"80",x"75",x"48",x"ed"),
  1897 => (x"97",x"6e",x"7e",x"70"),
  1898 => (x"4b",x"49",x"4b",x"bf"),
  1899 => (x"a3",x"c1",x"48",x"6e"),
  1900 => (x"11",x"81",x"6a",x"50"),
  1901 => (x"58",x"a6",x"cc",x"48"),
  1902 => (x"c4",x"02",x"ac",x"70"),
  1903 => (x"c0",x"48",x"6e",x"87"),
  1904 => (x"05",x"66",x"c8",x"50"),
  1905 => (x"f5",x"c2",x"87",x"c7"),
  1906 => (x"a5",x"c4",x"48",x"f1"),
  1907 => (x"c4",x"85",x"c1",x"78"),
  1908 => (x"ff",x"04",x"ad",x"b7"),
  1909 => (x"dc",x"c4",x"87",x"c0"),
  1910 => (x"fd",x"f5",x"c2",x"87"),
  1911 => (x"b7",x"c8",x"48",x"bf"),
  1912 => (x"87",x"d1",x"01",x"a8"),
  1913 => (x"cc",x"02",x"ac",x"ca"),
  1914 => (x"02",x"ac",x"cd",x"87"),
  1915 => (x"b7",x"c0",x"87",x"c7"),
  1916 => (x"f3",x"c0",x"03",x"ac"),
  1917 => (x"fd",x"f5",x"c2",x"87"),
  1918 => (x"b7",x"c8",x"4b",x"bf"),
  1919 => (x"87",x"d2",x"03",x"ab"),
  1920 => (x"49",x"c1",x"f6",x"c2"),
  1921 => (x"e0",x"c0",x"81",x"73"),
  1922 => (x"c8",x"83",x"c1",x"51"),
  1923 => (x"ff",x"04",x"ab",x"b7"),
  1924 => (x"f6",x"c2",x"87",x"ee"),
  1925 => (x"d2",x"c1",x"48",x"c9"),
  1926 => (x"50",x"cf",x"c1",x"50"),
  1927 => (x"c0",x"50",x"cd",x"c1"),
  1928 => (x"c3",x"80",x"e4",x"50"),
  1929 => (x"87",x"cd",x"c3",x"78"),
  1930 => (x"bf",x"fd",x"f5",x"c2"),
  1931 => (x"80",x"c1",x"48",x"49"),
  1932 => (x"58",x"c1",x"f6",x"c2"),
  1933 => (x"81",x"a0",x"c4",x"48"),
  1934 => (x"f8",x"c2",x"51",x"74"),
  1935 => (x"b7",x"f0",x"c0",x"87"),
  1936 => (x"87",x"da",x"04",x"ac"),
  1937 => (x"ac",x"b7",x"f9",x"c0"),
  1938 => (x"c2",x"87",x"d3",x"01"),
  1939 => (x"49",x"bf",x"f5",x"f5"),
  1940 => (x"4a",x"74",x"91",x"ca"),
  1941 => (x"c2",x"8a",x"f0",x"c0"),
  1942 => (x"72",x"48",x"f5",x"f5"),
  1943 => (x"ac",x"ca",x"78",x"a1"),
  1944 => (x"87",x"c6",x"c0",x"02"),
  1945 => (x"c2",x"05",x"ac",x"cd"),
  1946 => (x"f5",x"c2",x"87",x"cb"),
  1947 => (x"78",x"c3",x"48",x"f1"),
  1948 => (x"c0",x"87",x"c2",x"c2"),
  1949 => (x"04",x"ac",x"b7",x"f0"),
  1950 => (x"f9",x"c0",x"87",x"db"),
  1951 => (x"c0",x"01",x"ac",x"b7"),
  1952 => (x"f5",x"c2",x"87",x"d3"),
  1953 => (x"d0",x"49",x"bf",x"f9"),
  1954 => (x"c0",x"4a",x"74",x"91"),
  1955 => (x"f5",x"c2",x"8a",x"f0"),
  1956 => (x"a1",x"72",x"48",x"f9"),
  1957 => (x"b7",x"c1",x"c1",x"78"),
  1958 => (x"db",x"c0",x"04",x"ac"),
  1959 => (x"b7",x"c6",x"c1",x"87"),
  1960 => (x"d3",x"c0",x"01",x"ac"),
  1961 => (x"f9",x"f5",x"c2",x"87"),
  1962 => (x"91",x"d0",x"49",x"bf"),
  1963 => (x"f7",x"c0",x"4a",x"74"),
  1964 => (x"f9",x"f5",x"c2",x"8a"),
  1965 => (x"78",x"a1",x"72",x"48"),
  1966 => (x"c0",x"02",x"ac",x"ca"),
  1967 => (x"ac",x"cd",x"87",x"c6"),
  1968 => (x"87",x"f1",x"c0",x"05"),
  1969 => (x"48",x"f1",x"f5",x"c2"),
  1970 => (x"e8",x"c0",x"78",x"c3"),
  1971 => (x"ac",x"e2",x"c0",x"87"),
  1972 => (x"87",x"c9",x"c0",x"05"),
  1973 => (x"c0",x"48",x"a6",x"c4"),
  1974 => (x"d8",x"c0",x"78",x"fb"),
  1975 => (x"02",x"ac",x"ca",x"87"),
  1976 => (x"cd",x"87",x"c6",x"c0"),
  1977 => (x"c9",x"c0",x"05",x"ac"),
  1978 => (x"f1",x"f5",x"c2",x"87"),
  1979 => (x"c0",x"78",x"c3",x"48"),
  1980 => (x"a6",x"c8",x"87",x"c3"),
  1981 => (x"ac",x"b7",x"c0",x"5c"),
  1982 => (x"87",x"c4",x"c0",x"03"),
  1983 => (x"87",x"ca",x"c0",x"48"),
  1984 => (x"f9",x"02",x"66",x"c4"),
  1985 => (x"c3",x"48",x"87",x"c6"),
  1986 => (x"8e",x"f4",x"99",x"ff"),
  1987 => (x"43",x"87",x"cf",x"f8"),
  1988 => (x"3d",x"46",x"4e",x"4f"),
  1989 => (x"44",x"4f",x"4d",x"00"),
  1990 => (x"4d",x"41",x"4e",x"00"),
  1991 => (x"45",x"44",x"00",x"45"),
  1992 => (x"4c",x"55",x"41",x"46"),
  1993 => (x"00",x"30",x"3d",x"54"),
  1994 => (x"00",x"00",x"1f",x"0f"),
  1995 => (x"00",x"00",x"1f",x"15"),
  1996 => (x"00",x"00",x"1f",x"19"),
  1997 => (x"00",x"00",x"1f",x"1e"),
  1998 => (x"48",x"d0",x"ff",x"1e"),
  1999 => (x"71",x"78",x"c9",x"c8"),
  2000 => (x"08",x"d4",x"ff",x"48"),
  2001 => (x"1e",x"4f",x"26",x"78"),
  2002 => (x"eb",x"49",x"4a",x"71"),
  2003 => (x"48",x"d0",x"ff",x"87"),
  2004 => (x"4f",x"26",x"78",x"c8"),
  2005 => (x"71",x"1e",x"73",x"1e"),
  2006 => (x"d9",x"f6",x"c2",x"4b"),
  2007 => (x"87",x"c3",x"02",x"bf"),
  2008 => (x"ff",x"87",x"eb",x"c2"),
  2009 => (x"c9",x"c8",x"48",x"d0"),
  2010 => (x"c0",x"49",x"73",x"78"),
  2011 => (x"d4",x"ff",x"b1",x"e0"),
  2012 => (x"c2",x"78",x"71",x"48"),
  2013 => (x"c0",x"48",x"cd",x"f6"),
  2014 => (x"02",x"66",x"c8",x"78"),
  2015 => (x"ff",x"c3",x"87",x"c5"),
  2016 => (x"c0",x"87",x"c2",x"49"),
  2017 => (x"d5",x"f6",x"c2",x"49"),
  2018 => (x"02",x"66",x"cc",x"59"),
  2019 => (x"d5",x"c5",x"87",x"c6"),
  2020 => (x"87",x"c4",x"4a",x"d5"),
  2021 => (x"4a",x"ff",x"ff",x"cf"),
  2022 => (x"5a",x"d9",x"f6",x"c2"),
  2023 => (x"48",x"d9",x"f6",x"c2"),
  2024 => (x"87",x"c4",x"78",x"c1"),
  2025 => (x"4c",x"26",x"4d",x"26"),
  2026 => (x"4f",x"26",x"4b",x"26"),
  2027 => (x"5c",x"5b",x"5e",x"0e"),
  2028 => (x"4a",x"71",x"0e",x"5d"),
  2029 => (x"bf",x"d5",x"f6",x"c2"),
  2030 => (x"02",x"9a",x"72",x"4c"),
  2031 => (x"c8",x"49",x"87",x"cb"),
  2032 => (x"ca",x"fd",x"c1",x"91"),
  2033 => (x"c4",x"83",x"71",x"4b"),
  2034 => (x"ca",x"c1",x"c2",x"87"),
  2035 => (x"13",x"4d",x"c0",x"4b"),
  2036 => (x"c2",x"99",x"74",x"49"),
  2037 => (x"b9",x"bf",x"d1",x"f6"),
  2038 => (x"71",x"48",x"d4",x"ff"),
  2039 => (x"2c",x"b7",x"c1",x"78"),
  2040 => (x"ad",x"b7",x"c8",x"85"),
  2041 => (x"c2",x"87",x"e8",x"04"),
  2042 => (x"48",x"bf",x"cd",x"f6"),
  2043 => (x"f6",x"c2",x"80",x"c8"),
  2044 => (x"ef",x"fe",x"58",x"d1"),
  2045 => (x"1e",x"73",x"1e",x"87"),
  2046 => (x"4a",x"13",x"4b",x"71"),
  2047 => (x"87",x"cb",x"02",x"9a"),
  2048 => (x"e7",x"fe",x"49",x"72"),
  2049 => (x"9a",x"4a",x"13",x"87"),
  2050 => (x"fe",x"87",x"f5",x"05"),
  2051 => (x"c2",x"1e",x"87",x"da"),
  2052 => (x"49",x"bf",x"cd",x"f6"),
  2053 => (x"48",x"cd",x"f6",x"c2"),
  2054 => (x"c4",x"78",x"a1",x"c1"),
  2055 => (x"03",x"a9",x"b7",x"c0"),
  2056 => (x"d4",x"ff",x"87",x"db"),
  2057 => (x"d1",x"f6",x"c2",x"48"),
  2058 => (x"f6",x"c2",x"78",x"bf"),
  2059 => (x"c2",x"49",x"bf",x"cd"),
  2060 => (x"c1",x"48",x"cd",x"f6"),
  2061 => (x"c0",x"c4",x"78",x"a1"),
  2062 => (x"e5",x"04",x"a9",x"b7"),
  2063 => (x"48",x"d0",x"ff",x"87"),
  2064 => (x"f6",x"c2",x"78",x"c8"),
  2065 => (x"78",x"c0",x"48",x"d9"),
  2066 => (x"00",x"00",x"4f",x"26"),
  2067 => (x"00",x"00",x"00",x"00"),
  2068 => (x"00",x"00",x"00",x"00"),
  2069 => (x"00",x"5f",x"5f",x"00"),
  2070 => (x"03",x"00",x"00",x"00"),
  2071 => (x"03",x"03",x"00",x"03"),
  2072 => (x"7f",x"14",x"00",x"00"),
  2073 => (x"7f",x"7f",x"14",x"7f"),
  2074 => (x"24",x"00",x"00",x"14"),
  2075 => (x"3a",x"6b",x"6b",x"2e"),
  2076 => (x"6a",x"4c",x"00",x"12"),
  2077 => (x"56",x"6c",x"18",x"36"),
  2078 => (x"7e",x"30",x"00",x"32"),
  2079 => (x"3a",x"77",x"59",x"4f"),
  2080 => (x"00",x"00",x"40",x"68"),
  2081 => (x"00",x"03",x"07",x"04"),
  2082 => (x"00",x"00",x"00",x"00"),
  2083 => (x"41",x"63",x"3e",x"1c"),
  2084 => (x"00",x"00",x"00",x"00"),
  2085 => (x"1c",x"3e",x"63",x"41"),
  2086 => (x"2a",x"08",x"00",x"00"),
  2087 => (x"3e",x"1c",x"1c",x"3e"),
  2088 => (x"08",x"00",x"08",x"2a"),
  2089 => (x"08",x"3e",x"3e",x"08"),
  2090 => (x"00",x"00",x"00",x"08"),
  2091 => (x"00",x"60",x"e0",x"80"),
  2092 => (x"08",x"00",x"00",x"00"),
  2093 => (x"08",x"08",x"08",x"08"),
  2094 => (x"00",x"00",x"00",x"08"),
  2095 => (x"00",x"60",x"60",x"00"),
  2096 => (x"60",x"40",x"00",x"00"),
  2097 => (x"06",x"0c",x"18",x"30"),
  2098 => (x"3e",x"00",x"01",x"03"),
  2099 => (x"7f",x"4d",x"59",x"7f"),
  2100 => (x"04",x"00",x"00",x"3e"),
  2101 => (x"00",x"7f",x"7f",x"06"),
  2102 => (x"42",x"00",x"00",x"00"),
  2103 => (x"4f",x"59",x"71",x"63"),
  2104 => (x"22",x"00",x"00",x"46"),
  2105 => (x"7f",x"49",x"49",x"63"),
  2106 => (x"1c",x"18",x"00",x"36"),
  2107 => (x"7f",x"7f",x"13",x"16"),
  2108 => (x"27",x"00",x"00",x"10"),
  2109 => (x"7d",x"45",x"45",x"67"),
  2110 => (x"3c",x"00",x"00",x"39"),
  2111 => (x"79",x"49",x"4b",x"7e"),
  2112 => (x"01",x"00",x"00",x"30"),
  2113 => (x"0f",x"79",x"71",x"01"),
  2114 => (x"36",x"00",x"00",x"07"),
  2115 => (x"7f",x"49",x"49",x"7f"),
  2116 => (x"06",x"00",x"00",x"36"),
  2117 => (x"3f",x"69",x"49",x"4f"),
  2118 => (x"00",x"00",x"00",x"1e"),
  2119 => (x"00",x"66",x"66",x"00"),
  2120 => (x"00",x"00",x"00",x"00"),
  2121 => (x"00",x"66",x"e6",x"80"),
  2122 => (x"08",x"00",x"00",x"00"),
  2123 => (x"22",x"14",x"14",x"08"),
  2124 => (x"14",x"00",x"00",x"22"),
  2125 => (x"14",x"14",x"14",x"14"),
  2126 => (x"22",x"00",x"00",x"14"),
  2127 => (x"08",x"14",x"14",x"22"),
  2128 => (x"02",x"00",x"00",x"08"),
  2129 => (x"0f",x"59",x"51",x"03"),
  2130 => (x"7f",x"3e",x"00",x"06"),
  2131 => (x"1f",x"55",x"5d",x"41"),
  2132 => (x"7e",x"00",x"00",x"1e"),
  2133 => (x"7f",x"09",x"09",x"7f"),
  2134 => (x"7f",x"00",x"00",x"7e"),
  2135 => (x"7f",x"49",x"49",x"7f"),
  2136 => (x"1c",x"00",x"00",x"36"),
  2137 => (x"41",x"41",x"63",x"3e"),
  2138 => (x"7f",x"00",x"00",x"41"),
  2139 => (x"3e",x"63",x"41",x"7f"),
  2140 => (x"7f",x"00",x"00",x"1c"),
  2141 => (x"41",x"49",x"49",x"7f"),
  2142 => (x"7f",x"00",x"00",x"41"),
  2143 => (x"01",x"09",x"09",x"7f"),
  2144 => (x"3e",x"00",x"00",x"01"),
  2145 => (x"7b",x"49",x"41",x"7f"),
  2146 => (x"7f",x"00",x"00",x"7a"),
  2147 => (x"7f",x"08",x"08",x"7f"),
  2148 => (x"00",x"00",x"00",x"7f"),
  2149 => (x"41",x"7f",x"7f",x"41"),
  2150 => (x"20",x"00",x"00",x"00"),
  2151 => (x"7f",x"40",x"40",x"60"),
  2152 => (x"7f",x"7f",x"00",x"3f"),
  2153 => (x"63",x"36",x"1c",x"08"),
  2154 => (x"7f",x"00",x"00",x"41"),
  2155 => (x"40",x"40",x"40",x"7f"),
  2156 => (x"7f",x"7f",x"00",x"40"),
  2157 => (x"7f",x"06",x"0c",x"06"),
  2158 => (x"7f",x"7f",x"00",x"7f"),
  2159 => (x"7f",x"18",x"0c",x"06"),
  2160 => (x"3e",x"00",x"00",x"7f"),
  2161 => (x"7f",x"41",x"41",x"7f"),
  2162 => (x"7f",x"00",x"00",x"3e"),
  2163 => (x"0f",x"09",x"09",x"7f"),
  2164 => (x"7f",x"3e",x"00",x"06"),
  2165 => (x"7e",x"7f",x"61",x"41"),
  2166 => (x"7f",x"00",x"00",x"40"),
  2167 => (x"7f",x"19",x"09",x"7f"),
  2168 => (x"26",x"00",x"00",x"66"),
  2169 => (x"7b",x"59",x"4d",x"6f"),
  2170 => (x"01",x"00",x"00",x"32"),
  2171 => (x"01",x"7f",x"7f",x"01"),
  2172 => (x"3f",x"00",x"00",x"01"),
  2173 => (x"7f",x"40",x"40",x"7f"),
  2174 => (x"0f",x"00",x"00",x"3f"),
  2175 => (x"3f",x"70",x"70",x"3f"),
  2176 => (x"7f",x"7f",x"00",x"0f"),
  2177 => (x"7f",x"30",x"18",x"30"),
  2178 => (x"63",x"41",x"00",x"7f"),
  2179 => (x"36",x"1c",x"1c",x"36"),
  2180 => (x"03",x"01",x"41",x"63"),
  2181 => (x"06",x"7c",x"7c",x"06"),
  2182 => (x"71",x"61",x"01",x"03"),
  2183 => (x"43",x"47",x"4d",x"59"),
  2184 => (x"00",x"00",x"00",x"41"),
  2185 => (x"41",x"41",x"7f",x"7f"),
  2186 => (x"03",x"01",x"00",x"00"),
  2187 => (x"30",x"18",x"0c",x"06"),
  2188 => (x"00",x"00",x"40",x"60"),
  2189 => (x"7f",x"7f",x"41",x"41"),
  2190 => (x"0c",x"08",x"00",x"00"),
  2191 => (x"0c",x"06",x"03",x"06"),
  2192 => (x"80",x"80",x"00",x"08"),
  2193 => (x"80",x"80",x"80",x"80"),
  2194 => (x"00",x"00",x"00",x"80"),
  2195 => (x"04",x"07",x"03",x"00"),
  2196 => (x"20",x"00",x"00",x"00"),
  2197 => (x"7c",x"54",x"54",x"74"),
  2198 => (x"7f",x"00",x"00",x"78"),
  2199 => (x"7c",x"44",x"44",x"7f"),
  2200 => (x"38",x"00",x"00",x"38"),
  2201 => (x"44",x"44",x"44",x"7c"),
  2202 => (x"38",x"00",x"00",x"00"),
  2203 => (x"7f",x"44",x"44",x"7c"),
  2204 => (x"38",x"00",x"00",x"7f"),
  2205 => (x"5c",x"54",x"54",x"7c"),
  2206 => (x"04",x"00",x"00",x"18"),
  2207 => (x"05",x"05",x"7f",x"7e"),
  2208 => (x"18",x"00",x"00",x"00"),
  2209 => (x"fc",x"a4",x"a4",x"bc"),
  2210 => (x"7f",x"00",x"00",x"7c"),
  2211 => (x"7c",x"04",x"04",x"7f"),
  2212 => (x"00",x"00",x"00",x"78"),
  2213 => (x"40",x"7d",x"3d",x"00"),
  2214 => (x"80",x"00",x"00",x"00"),
  2215 => (x"7d",x"fd",x"80",x"80"),
  2216 => (x"7f",x"00",x"00",x"00"),
  2217 => (x"6c",x"38",x"10",x"7f"),
  2218 => (x"00",x"00",x"00",x"44"),
  2219 => (x"40",x"7f",x"3f",x"00"),
  2220 => (x"7c",x"7c",x"00",x"00"),
  2221 => (x"7c",x"0c",x"18",x"0c"),
  2222 => (x"7c",x"00",x"00",x"78"),
  2223 => (x"7c",x"04",x"04",x"7c"),
  2224 => (x"38",x"00",x"00",x"78"),
  2225 => (x"7c",x"44",x"44",x"7c"),
  2226 => (x"fc",x"00",x"00",x"38"),
  2227 => (x"3c",x"24",x"24",x"fc"),
  2228 => (x"18",x"00",x"00",x"18"),
  2229 => (x"fc",x"24",x"24",x"3c"),
  2230 => (x"7c",x"00",x"00",x"fc"),
  2231 => (x"0c",x"04",x"04",x"7c"),
  2232 => (x"48",x"00",x"00",x"08"),
  2233 => (x"74",x"54",x"54",x"5c"),
  2234 => (x"04",x"00",x"00",x"20"),
  2235 => (x"44",x"44",x"7f",x"3f"),
  2236 => (x"3c",x"00",x"00",x"00"),
  2237 => (x"7c",x"40",x"40",x"7c"),
  2238 => (x"1c",x"00",x"00",x"7c"),
  2239 => (x"3c",x"60",x"60",x"3c"),
  2240 => (x"7c",x"3c",x"00",x"1c"),
  2241 => (x"7c",x"60",x"30",x"60"),
  2242 => (x"6c",x"44",x"00",x"3c"),
  2243 => (x"6c",x"38",x"10",x"38"),
  2244 => (x"1c",x"00",x"00",x"44"),
  2245 => (x"3c",x"60",x"e0",x"bc"),
  2246 => (x"44",x"00",x"00",x"1c"),
  2247 => (x"4c",x"5c",x"74",x"64"),
  2248 => (x"08",x"00",x"00",x"44"),
  2249 => (x"41",x"77",x"3e",x"08"),
  2250 => (x"00",x"00",x"00",x"41"),
  2251 => (x"00",x"7f",x"7f",x"00"),
  2252 => (x"41",x"00",x"00",x"00"),
  2253 => (x"08",x"3e",x"77",x"41"),
  2254 => (x"01",x"02",x"00",x"08"),
  2255 => (x"02",x"02",x"03",x"01"),
  2256 => (x"7f",x"7f",x"00",x"01"),
  2257 => (x"7f",x"7f",x"7f",x"7f"),
  2258 => (x"08",x"08",x"00",x"7f"),
  2259 => (x"3e",x"3e",x"1c",x"1c"),
  2260 => (x"7f",x"7f",x"7f",x"7f"),
  2261 => (x"1c",x"1c",x"3e",x"3e"),
  2262 => (x"10",x"00",x"08",x"08"),
  2263 => (x"18",x"7c",x"7c",x"18"),
  2264 => (x"10",x"00",x"00",x"10"),
  2265 => (x"30",x"7c",x"7c",x"30"),
  2266 => (x"30",x"10",x"00",x"10"),
  2267 => (x"1e",x"78",x"60",x"60"),
  2268 => (x"66",x"42",x"00",x"06"),
  2269 => (x"66",x"3c",x"18",x"3c"),
  2270 => (x"38",x"78",x"00",x"42"),
  2271 => (x"6c",x"c6",x"c2",x"6a"),
  2272 => (x"00",x"60",x"00",x"38"),
  2273 => (x"00",x"00",x"60",x"00"),
  2274 => (x"5e",x"0e",x"00",x"60"),
  2275 => (x"0e",x"5d",x"5c",x"5b"),
  2276 => (x"c2",x"4c",x"71",x"1e"),
  2277 => (x"4d",x"bf",x"ea",x"f6"),
  2278 => (x"1e",x"c0",x"4b",x"c0"),
  2279 => (x"c7",x"02",x"ab",x"74"),
  2280 => (x"48",x"a6",x"c4",x"87"),
  2281 => (x"87",x"c5",x"78",x"c0"),
  2282 => (x"c1",x"48",x"a6",x"c4"),
  2283 => (x"1e",x"66",x"c4",x"78"),
  2284 => (x"df",x"ee",x"49",x"73"),
  2285 => (x"c0",x"86",x"c8",x"87"),
  2286 => (x"ef",x"ef",x"49",x"e0"),
  2287 => (x"4a",x"a5",x"c4",x"87"),
  2288 => (x"f0",x"f0",x"49",x"6a"),
  2289 => (x"87",x"c6",x"f1",x"87"),
  2290 => (x"83",x"c1",x"85",x"cb"),
  2291 => (x"04",x"ab",x"b7",x"c8"),
  2292 => (x"26",x"87",x"c7",x"ff"),
  2293 => (x"4c",x"26",x"4d",x"26"),
  2294 => (x"4f",x"26",x"4b",x"26"),
  2295 => (x"c2",x"4a",x"71",x"1e"),
  2296 => (x"c2",x"5a",x"ee",x"f6"),
  2297 => (x"c7",x"48",x"ee",x"f6"),
  2298 => (x"dd",x"fe",x"49",x"78"),
  2299 => (x"1e",x"4f",x"26",x"87"),
  2300 => (x"4a",x"71",x"1e",x"73"),
  2301 => (x"03",x"aa",x"b7",x"c0"),
  2302 => (x"dd",x"c2",x"87",x"d3"),
  2303 => (x"c4",x"05",x"bf",x"cf"),
  2304 => (x"c2",x"4b",x"c1",x"87"),
  2305 => (x"c2",x"4b",x"c0",x"87"),
  2306 => (x"c4",x"5b",x"d3",x"dd"),
  2307 => (x"d3",x"dd",x"c2",x"87"),
  2308 => (x"cf",x"dd",x"c2",x"5a"),
  2309 => (x"9a",x"c1",x"4a",x"bf"),
  2310 => (x"49",x"a2",x"c0",x"c1"),
  2311 => (x"fc",x"87",x"e8",x"ec"),
  2312 => (x"cf",x"dd",x"c2",x"48"),
  2313 => (x"ef",x"fe",x"78",x"bf"),
  2314 => (x"4a",x"71",x"1e",x"87"),
  2315 => (x"72",x"1e",x"66",x"c4"),
  2316 => (x"da",x"df",x"ff",x"49"),
  2317 => (x"4f",x"26",x"26",x"87"),
  2318 => (x"cf",x"dd",x"c2",x"1e"),
  2319 => (x"dc",x"ff",x"49",x"bf"),
  2320 => (x"f6",x"c2",x"87",x"c2"),
  2321 => (x"bf",x"e8",x"48",x"e2"),
  2322 => (x"de",x"f6",x"c2",x"78"),
  2323 => (x"78",x"bf",x"ec",x"48"),
  2324 => (x"bf",x"e2",x"f6",x"c2"),
  2325 => (x"ff",x"c3",x"49",x"4a"),
  2326 => (x"2a",x"b7",x"c8",x"99"),
  2327 => (x"b0",x"71",x"48",x"72"),
  2328 => (x"58",x"ea",x"f6",x"c2"),
  2329 => (x"5e",x"0e",x"4f",x"26"),
  2330 => (x"0e",x"5d",x"5c",x"5b"),
  2331 => (x"c7",x"ff",x"4b",x"71"),
  2332 => (x"dd",x"f6",x"c2",x"87"),
  2333 => (x"73",x"50",x"c0",x"48"),
  2334 => (x"e7",x"db",x"ff",x"49"),
  2335 => (x"4c",x"49",x"70",x"87"),
  2336 => (x"ee",x"cb",x"9c",x"c2"),
  2337 => (x"87",x"cf",x"cb",x"49"),
  2338 => (x"c2",x"4d",x"49",x"70"),
  2339 => (x"bf",x"97",x"dd",x"f6"),
  2340 => (x"87",x"e4",x"c1",x"05"),
  2341 => (x"c2",x"49",x"66",x"d0"),
  2342 => (x"99",x"bf",x"e6",x"f6"),
  2343 => (x"d4",x"87",x"d7",x"05"),
  2344 => (x"f6",x"c2",x"49",x"66"),
  2345 => (x"05",x"99",x"bf",x"de"),
  2346 => (x"49",x"73",x"87",x"cc"),
  2347 => (x"87",x"f4",x"da",x"ff"),
  2348 => (x"c1",x"02",x"98",x"70"),
  2349 => (x"4c",x"c1",x"87",x"c2"),
  2350 => (x"75",x"87",x"fd",x"fd"),
  2351 => (x"87",x"e3",x"ca",x"49"),
  2352 => (x"c6",x"02",x"98",x"70"),
  2353 => (x"dd",x"f6",x"c2",x"87"),
  2354 => (x"c2",x"50",x"c1",x"48"),
  2355 => (x"bf",x"97",x"dd",x"f6"),
  2356 => (x"87",x"e4",x"c0",x"05"),
  2357 => (x"bf",x"e6",x"f6",x"c2"),
  2358 => (x"99",x"66",x"d0",x"49"),
  2359 => (x"87",x"d6",x"ff",x"05"),
  2360 => (x"bf",x"de",x"f6",x"c2"),
  2361 => (x"99",x"66",x"d4",x"49"),
  2362 => (x"87",x"ca",x"ff",x"05"),
  2363 => (x"d9",x"ff",x"49",x"73"),
  2364 => (x"98",x"70",x"87",x"f2"),
  2365 => (x"87",x"fe",x"fe",x"05"),
  2366 => (x"d7",x"fb",x"48",x"74"),
  2367 => (x"5b",x"5e",x"0e",x"87"),
  2368 => (x"f4",x"0e",x"5d",x"5c"),
  2369 => (x"4c",x"4d",x"c0",x"86"),
  2370 => (x"c4",x"7e",x"bf",x"ec"),
  2371 => (x"f6",x"c2",x"48",x"a6"),
  2372 => (x"c1",x"78",x"bf",x"ea"),
  2373 => (x"c7",x"1e",x"c0",x"1e"),
  2374 => (x"87",x"ca",x"fd",x"49"),
  2375 => (x"98",x"70",x"86",x"c8"),
  2376 => (x"ff",x"87",x"ce",x"02"),
  2377 => (x"87",x"c7",x"fb",x"49"),
  2378 => (x"ff",x"49",x"da",x"c1"),
  2379 => (x"c1",x"87",x"f5",x"d8"),
  2380 => (x"dd",x"f6",x"c2",x"4d"),
  2381 => (x"c3",x"02",x"bf",x"97"),
  2382 => (x"87",x"f9",x"cd",x"87"),
  2383 => (x"bf",x"e2",x"f6",x"c2"),
  2384 => (x"cf",x"dd",x"c2",x"4b"),
  2385 => (x"eb",x"c0",x"05",x"bf"),
  2386 => (x"49",x"fd",x"c3",x"87"),
  2387 => (x"87",x"d4",x"d8",x"ff"),
  2388 => (x"ff",x"49",x"fa",x"c3"),
  2389 => (x"73",x"87",x"cd",x"d8"),
  2390 => (x"99",x"ff",x"c3",x"49"),
  2391 => (x"49",x"c0",x"1e",x"71"),
  2392 => (x"73",x"87",x"c6",x"fb"),
  2393 => (x"29",x"b7",x"c8",x"49"),
  2394 => (x"49",x"c1",x"1e",x"71"),
  2395 => (x"c8",x"87",x"fa",x"fa"),
  2396 => (x"87",x"c1",x"c6",x"86"),
  2397 => (x"bf",x"e6",x"f6",x"c2"),
  2398 => (x"dd",x"02",x"9b",x"4b"),
  2399 => (x"cb",x"dd",x"c2",x"87"),
  2400 => (x"de",x"c7",x"49",x"bf"),
  2401 => (x"05",x"98",x"70",x"87"),
  2402 => (x"4b",x"c0",x"87",x"c4"),
  2403 => (x"e0",x"c2",x"87",x"d2"),
  2404 => (x"87",x"c3",x"c7",x"49"),
  2405 => (x"58",x"cf",x"dd",x"c2"),
  2406 => (x"dd",x"c2",x"87",x"c6"),
  2407 => (x"78",x"c0",x"48",x"cb"),
  2408 => (x"99",x"c2",x"49",x"73"),
  2409 => (x"c3",x"87",x"ce",x"05"),
  2410 => (x"d6",x"ff",x"49",x"eb"),
  2411 => (x"49",x"70",x"87",x"f6"),
  2412 => (x"c2",x"02",x"99",x"c2"),
  2413 => (x"73",x"4c",x"fb",x"87"),
  2414 => (x"05",x"99",x"c1",x"49"),
  2415 => (x"f4",x"c3",x"87",x"ce"),
  2416 => (x"df",x"d6",x"ff",x"49"),
  2417 => (x"c2",x"49",x"70",x"87"),
  2418 => (x"87",x"c2",x"02",x"99"),
  2419 => (x"49",x"73",x"4c",x"fa"),
  2420 => (x"ce",x"05",x"99",x"c8"),
  2421 => (x"49",x"f5",x"c3",x"87"),
  2422 => (x"87",x"c8",x"d6",x"ff"),
  2423 => (x"99",x"c2",x"49",x"70"),
  2424 => (x"c2",x"87",x"d5",x"02"),
  2425 => (x"02",x"bf",x"ee",x"f6"),
  2426 => (x"c1",x"48",x"87",x"ca"),
  2427 => (x"f2",x"f6",x"c2",x"88"),
  2428 => (x"87",x"c2",x"c0",x"58"),
  2429 => (x"4d",x"c1",x"4c",x"ff"),
  2430 => (x"99",x"c4",x"49",x"73"),
  2431 => (x"c3",x"87",x"ce",x"05"),
  2432 => (x"d5",x"ff",x"49",x"f2"),
  2433 => (x"49",x"70",x"87",x"de"),
  2434 => (x"dc",x"02",x"99",x"c2"),
  2435 => (x"ee",x"f6",x"c2",x"87"),
  2436 => (x"c7",x"48",x"7e",x"bf"),
  2437 => (x"c0",x"03",x"a8",x"b7"),
  2438 => (x"48",x"6e",x"87",x"cb"),
  2439 => (x"f6",x"c2",x"80",x"c1"),
  2440 => (x"c2",x"c0",x"58",x"f2"),
  2441 => (x"c1",x"4c",x"fe",x"87"),
  2442 => (x"49",x"fd",x"c3",x"4d"),
  2443 => (x"87",x"f4",x"d4",x"ff"),
  2444 => (x"99",x"c2",x"49",x"70"),
  2445 => (x"87",x"d5",x"c0",x"02"),
  2446 => (x"bf",x"ee",x"f6",x"c2"),
  2447 => (x"87",x"c9",x"c0",x"02"),
  2448 => (x"48",x"ee",x"f6",x"c2"),
  2449 => (x"c2",x"c0",x"78",x"c0"),
  2450 => (x"c1",x"4c",x"fd",x"87"),
  2451 => (x"49",x"fa",x"c3",x"4d"),
  2452 => (x"87",x"d0",x"d4",x"ff"),
  2453 => (x"99",x"c2",x"49",x"70"),
  2454 => (x"87",x"d9",x"c0",x"02"),
  2455 => (x"bf",x"ee",x"f6",x"c2"),
  2456 => (x"a8",x"b7",x"c7",x"48"),
  2457 => (x"87",x"c9",x"c0",x"03"),
  2458 => (x"48",x"ee",x"f6",x"c2"),
  2459 => (x"c2",x"c0",x"78",x"c7"),
  2460 => (x"c1",x"4c",x"fc",x"87"),
  2461 => (x"ac",x"b7",x"c0",x"4d"),
  2462 => (x"87",x"d1",x"c0",x"03"),
  2463 => (x"c1",x"4a",x"66",x"c4"),
  2464 => (x"02",x"6a",x"82",x"d8"),
  2465 => (x"6a",x"87",x"c6",x"c0"),
  2466 => (x"73",x"49",x"74",x"4b"),
  2467 => (x"c3",x"1e",x"c0",x"0f"),
  2468 => (x"da",x"c1",x"1e",x"f0"),
  2469 => (x"87",x"ce",x"f7",x"49"),
  2470 => (x"98",x"70",x"86",x"c8"),
  2471 => (x"87",x"e2",x"c0",x"02"),
  2472 => (x"c2",x"48",x"a6",x"c8"),
  2473 => (x"78",x"bf",x"ee",x"f6"),
  2474 => (x"cb",x"49",x"66",x"c8"),
  2475 => (x"48",x"66",x"c4",x"91"),
  2476 => (x"7e",x"70",x"80",x"71"),
  2477 => (x"c0",x"02",x"bf",x"6e"),
  2478 => (x"bf",x"6e",x"87",x"c8"),
  2479 => (x"49",x"66",x"c8",x"4b"),
  2480 => (x"9d",x"75",x"0f",x"73"),
  2481 => (x"87",x"c8",x"c0",x"02"),
  2482 => (x"bf",x"ee",x"f6",x"c2"),
  2483 => (x"87",x"fa",x"f2",x"49"),
  2484 => (x"bf",x"d3",x"dd",x"c2"),
  2485 => (x"87",x"dd",x"c0",x"02"),
  2486 => (x"87",x"c7",x"c2",x"49"),
  2487 => (x"c0",x"02",x"98",x"70"),
  2488 => (x"f6",x"c2",x"87",x"d3"),
  2489 => (x"f2",x"49",x"bf",x"ee"),
  2490 => (x"49",x"c0",x"87",x"e0"),
  2491 => (x"c2",x"87",x"c0",x"f4"),
  2492 => (x"c0",x"48",x"d3",x"dd"),
  2493 => (x"f3",x"8e",x"f4",x"78"),
  2494 => (x"5e",x"0e",x"87",x"da"),
  2495 => (x"0e",x"5d",x"5c",x"5b"),
  2496 => (x"c2",x"4c",x"71",x"1e"),
  2497 => (x"49",x"bf",x"ea",x"f6"),
  2498 => (x"4d",x"a1",x"cd",x"c1"),
  2499 => (x"69",x"81",x"d1",x"c1"),
  2500 => (x"02",x"9c",x"74",x"7e"),
  2501 => (x"a5",x"c4",x"87",x"cf"),
  2502 => (x"c2",x"7b",x"74",x"4b"),
  2503 => (x"49",x"bf",x"ea",x"f6"),
  2504 => (x"6e",x"87",x"f9",x"f2"),
  2505 => (x"05",x"9c",x"74",x"7b"),
  2506 => (x"4b",x"c0",x"87",x"c4"),
  2507 => (x"4b",x"c1",x"87",x"c2"),
  2508 => (x"fa",x"f2",x"49",x"73"),
  2509 => (x"02",x"66",x"d4",x"87"),
  2510 => (x"da",x"49",x"87",x"c7"),
  2511 => (x"c2",x"4a",x"70",x"87"),
  2512 => (x"c2",x"4a",x"c0",x"87"),
  2513 => (x"26",x"5a",x"d7",x"dd"),
  2514 => (x"00",x"87",x"c9",x"f2"),
  2515 => (x"00",x"00",x"00",x"00"),
  2516 => (x"00",x"00",x"00",x"00"),
  2517 => (x"1e",x"00",x"00",x"00"),
  2518 => (x"c8",x"ff",x"4a",x"71"),
  2519 => (x"a1",x"72",x"49",x"bf"),
  2520 => (x"1e",x"4f",x"26",x"48"),
  2521 => (x"89",x"bf",x"c8",x"ff"),
  2522 => (x"c0",x"c0",x"c0",x"fe"),
  2523 => (x"01",x"a9",x"c0",x"c0"),
  2524 => (x"4a",x"c0",x"87",x"c4"),
  2525 => (x"4a",x"c1",x"87",x"c2"),
  2526 => (x"4f",x"26",x"48",x"72"),
  2527 => (x"5c",x"5b",x"5e",x"0e"),
  2528 => (x"71",x"1e",x"0e",x"5d"),
  2529 => (x"4b",x"d4",x"ff",x"4d"),
  2530 => (x"f6",x"c2",x"1e",x"75"),
  2531 => (x"c1",x"fe",x"49",x"f2"),
  2532 => (x"86",x"c4",x"87",x"d0"),
  2533 => (x"02",x"6e",x"7e",x"70"),
  2534 => (x"c2",x"87",x"ff",x"c3"),
  2535 => (x"4c",x"bf",x"fa",x"f6"),
  2536 => (x"da",x"fe",x"49",x"75"),
  2537 => (x"a8",x"de",x"87",x"fe"),
  2538 => (x"87",x"eb",x"c0",x"05"),
  2539 => (x"d3",x"ff",x"49",x"75"),
  2540 => (x"98",x"70",x"87",x"ec"),
  2541 => (x"c2",x"87",x"db",x"02"),
  2542 => (x"1e",x"bf",x"f5",x"f5"),
  2543 => (x"ff",x"49",x"e1",x"c0"),
  2544 => (x"c4",x"87",x"f7",x"d0"),
  2545 => (x"f4",x"e2",x"c2",x"86"),
  2546 => (x"c2",x"50",x"c0",x"48"),
  2547 => (x"fe",x"49",x"c1",x"f6"),
  2548 => (x"48",x"c1",x"87",x"ea"),
  2549 => (x"ff",x"87",x"c5",x"c3"),
  2550 => (x"c5",x"c8",x"48",x"d0"),
  2551 => (x"7b",x"d6",x"c1",x"78"),
  2552 => (x"97",x"6e",x"4a",x"c0"),
  2553 => (x"48",x"6e",x"7b",x"bf"),
  2554 => (x"7e",x"70",x"80",x"c1"),
  2555 => (x"e0",x"c0",x"82",x"c1"),
  2556 => (x"ff",x"04",x"aa",x"b7"),
  2557 => (x"d0",x"ff",x"87",x"ec"),
  2558 => (x"c8",x"78",x"c4",x"48"),
  2559 => (x"d3",x"c1",x"78",x"c5"),
  2560 => (x"c4",x"7b",x"c1",x"7b"),
  2561 => (x"02",x"9c",x"74",x"78"),
  2562 => (x"c2",x"87",x"fd",x"c1"),
  2563 => (x"c8",x"7e",x"ee",x"e4"),
  2564 => (x"c0",x"8c",x"4d",x"c0"),
  2565 => (x"c6",x"03",x"ac",x"b7"),
  2566 => (x"a4",x"c0",x"c8",x"87"),
  2567 => (x"c2",x"4c",x"c0",x"4d"),
  2568 => (x"bf",x"97",x"df",x"f1"),
  2569 => (x"02",x"99",x"d0",x"49"),
  2570 => (x"1e",x"c0",x"87",x"d2"),
  2571 => (x"49",x"f2",x"f6",x"c2"),
  2572 => (x"87",x"ca",x"c2",x"fe"),
  2573 => (x"49",x"70",x"86",x"c4"),
  2574 => (x"87",x"ef",x"c0",x"4a"),
  2575 => (x"1e",x"ee",x"e4",x"c2"),
  2576 => (x"49",x"f2",x"f6",x"c2"),
  2577 => (x"87",x"f6",x"c1",x"fe"),
  2578 => (x"49",x"70",x"86",x"c4"),
  2579 => (x"48",x"d0",x"ff",x"4a"),
  2580 => (x"c1",x"78",x"c5",x"c8"),
  2581 => (x"97",x"6e",x"7b",x"d4"),
  2582 => (x"48",x"6e",x"7b",x"bf"),
  2583 => (x"7e",x"70",x"80",x"c1"),
  2584 => (x"ff",x"05",x"8d",x"c1"),
  2585 => (x"d0",x"ff",x"87",x"f0"),
  2586 => (x"72",x"78",x"c4",x"48"),
  2587 => (x"c5",x"c0",x"05",x"9a"),
  2588 => (x"c0",x"48",x"c0",x"87"),
  2589 => (x"1e",x"c1",x"87",x"e6"),
  2590 => (x"49",x"f2",x"f6",x"c2"),
  2591 => (x"87",x"dd",x"ff",x"fd"),
  2592 => (x"9c",x"74",x"86",x"c4"),
  2593 => (x"87",x"c3",x"fe",x"05"),
  2594 => (x"c8",x"48",x"d0",x"ff"),
  2595 => (x"d3",x"c1",x"78",x"c5"),
  2596 => (x"c4",x"7b",x"c0",x"7b"),
  2597 => (x"c0",x"48",x"c1",x"78"),
  2598 => (x"48",x"c0",x"87",x"c2"),
  2599 => (x"26",x"4d",x"26",x"26"),
  2600 => (x"26",x"4b",x"26",x"4c"),
  2601 => (x"4a",x"71",x"1e",x"4f"),
  2602 => (x"c5",x"05",x"66",x"c4"),
  2603 => (x"fb",x"49",x"72",x"87"),
  2604 => (x"4f",x"26",x"87",x"ca"),
  2605 => (x"e4",x"c2",x"1e",x"00"),
  2606 => (x"c1",x"49",x"bf",x"c3"),
  2607 => (x"c7",x"e4",x"c2",x"b9"),
  2608 => (x"48",x"d4",x"ff",x"59"),
  2609 => (x"ff",x"78",x"ff",x"c3"),
  2610 => (x"e1",x"c8",x"48",x"d0"),
  2611 => (x"48",x"d4",x"ff",x"78"),
  2612 => (x"31",x"c4",x"78",x"c1"),
  2613 => (x"d0",x"ff",x"78",x"71"),
  2614 => (x"78",x"e0",x"c0",x"48"),
  2615 => (x"c2",x"1e",x"4f",x"26"),
  2616 => (x"c2",x"1e",x"f7",x"e3"),
  2617 => (x"fd",x"49",x"f2",x"f6"),
  2618 => (x"c4",x"87",x"f7",x"fb"),
  2619 => (x"02",x"98",x"70",x"86"),
  2620 => (x"c0",x"ff",x"87",x"c3"),
  2621 => (x"31",x"4f",x"26",x"87"),
  2622 => (x"5a",x"48",x"4b",x"35"),
  2623 => (x"43",x"20",x"20",x"20"),
  2624 => (x"00",x"00",x"47",x"46"),
  2625 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

