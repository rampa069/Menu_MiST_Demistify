library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c8f7c287",
    12 => x"86c0c64e",
    13 => x"49c8f7c2",
    14 => x"48c8e4c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087e1e0",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"ff1e4f26",
    53 => x"ffc348d4",
    54 => x"c4516878",
    55 => x"88c14866",
    56 => x"7058a6c8",
    57 => x"87eb0598",
    58 => x"731e4f26",
    59 => x"4bd4ff1e",
    60 => x"6b7bffc3",
    61 => x"7bffc34a",
    62 => x"32c8496b",
    63 => x"ffc3b172",
    64 => x"c84a6b7b",
    65 => x"c3b27131",
    66 => x"496b7bff",
    67 => x"b17232c8",
    68 => x"87c44871",
    69 => x"4c264d26",
    70 => x"4f264b26",
    71 => x"5c5b5e0e",
    72 => x"4a710e5d",
    73 => x"724cd4ff",
    74 => x"99ffc349",
    75 => x"e4c27c71",
    76 => x"c805bfc8",
    77 => x"4866d087",
    78 => x"a6d430c9",
    79 => x"4966d058",
    80 => x"ffc329d8",
    81 => x"d07c7199",
    82 => x"29d04966",
    83 => x"7199ffc3",
    84 => x"4966d07c",
    85 => x"ffc329c8",
    86 => x"d07c7199",
    87 => x"ffc34966",
    88 => x"727c7199",
    89 => x"c329d049",
    90 => x"7c7199ff",
    91 => x"f0c94b6c",
    92 => x"ffc34dff",
    93 => x"87d005ab",
    94 => x"6c7cffc3",
    95 => x"028dc14b",
    96 => x"ffc387c6",
    97 => x"87f002ab",
    98 => x"c7fe4873",
    99 => x"49c01e87",
   100 => x"c348d4ff",
   101 => x"81c178ff",
   102 => x"a9b7c8c3",
   103 => x"2687f104",
   104 => x"1e731e4f",
   105 => x"f8c487e7",
   106 => x"1ec04bdf",
   107 => x"c1f0ffc0",
   108 => x"e7fd49f7",
   109 => x"c186c487",
   110 => x"eac005a8",
   111 => x"48d4ff87",
   112 => x"c178ffc3",
   113 => x"c0c0c0c0",
   114 => x"e1c01ec0",
   115 => x"49e9c1f0",
   116 => x"c487c9fd",
   117 => x"05987086",
   118 => x"d4ff87ca",
   119 => x"78ffc348",
   120 => x"87cb48c1",
   121 => x"c187e6fe",
   122 => x"fdfe058b",
   123 => x"fc48c087",
   124 => x"731e87e6",
   125 => x"48d4ff1e",
   126 => x"d378ffc3",
   127 => x"c01ec04b",
   128 => x"c1c1f0ff",
   129 => x"87d4fc49",
   130 => x"987086c4",
   131 => x"ff87ca05",
   132 => x"ffc348d4",
   133 => x"cb48c178",
   134 => x"87f1fd87",
   135 => x"ff058bc1",
   136 => x"48c087db",
   137 => x"0e87f1fb",
   138 => x"0e5c5b5e",
   139 => x"fd4cd4ff",
   140 => x"eac687db",
   141 => x"f0e1c01e",
   142 => x"fb49c8c1",
   143 => x"86c487de",
   144 => x"c802a8c1",
   145 => x"87eafe87",
   146 => x"e2c148c0",
   147 => x"87dafa87",
   148 => x"ffcf4970",
   149 => x"eac699ff",
   150 => x"87c802a9",
   151 => x"c087d3fe",
   152 => x"87cbc148",
   153 => x"c07cffc3",
   154 => x"f4fc4bf1",
   155 => x"02987087",
   156 => x"c087ebc0",
   157 => x"f0ffc01e",
   158 => x"fa49fac1",
   159 => x"86c487de",
   160 => x"d9059870",
   161 => x"7cffc387",
   162 => x"ffc3496c",
   163 => x"7c7c7c7c",
   164 => x"0299c0c1",
   165 => x"48c187c4",
   166 => x"48c087d5",
   167 => x"abc287d1",
   168 => x"c087c405",
   169 => x"c187c848",
   170 => x"fdfe058b",
   171 => x"f948c087",
   172 => x"731e87e4",
   173 => x"c8e4c21e",
   174 => x"c778c148",
   175 => x"48d0ff4b",
   176 => x"c8fb78c2",
   177 => x"48d0ff87",
   178 => x"1ec078c3",
   179 => x"c1d0e5c0",
   180 => x"c7f949c0",
   181 => x"c186c487",
   182 => x"87c105a8",
   183 => x"05abc24b",
   184 => x"48c087c5",
   185 => x"c187f9c0",
   186 => x"d0ff058b",
   187 => x"87f7fc87",
   188 => x"58cce4c2",
   189 => x"cd059870",
   190 => x"c01ec187",
   191 => x"d0c1f0ff",
   192 => x"87d8f849",
   193 => x"d4ff86c4",
   194 => x"78ffc348",
   195 => x"c287fec2",
   196 => x"ff58d0e4",
   197 => x"78c248d0",
   198 => x"c348d4ff",
   199 => x"48c178ff",
   200 => x"1e87f5f7",
   201 => x"ff4ad4ff",
   202 => x"d1c448d0",
   203 => x"7affc378",
   204 => x"f80589c1",
   205 => x"1e4f2687",
   206 => x"4b711e73",
   207 => x"dfcdeec5",
   208 => x"48d4ff4a",
   209 => x"6878ffc3",
   210 => x"a8fec348",
   211 => x"c187c502",
   212 => x"87ed058a",
   213 => x"c5059a72",
   214 => x"c048c087",
   215 => x"9b7387ea",
   216 => x"c887cc02",
   217 => x"49731e66",
   218 => x"c487e7f5",
   219 => x"c887c686",
   220 => x"eefe4966",
   221 => x"48d4ff87",
   222 => x"7878ffc3",
   223 => x"c5059b73",
   224 => x"48d0ff87",
   225 => x"48c178d0",
   226 => x"1e87cdf6",
   227 => x"4a711e73",
   228 => x"d4ff4bc0",
   229 => x"78ffc348",
   230 => x"c448d0ff",
   231 => x"d4ff78c3",
   232 => x"78ffc348",
   233 => x"ffc01e72",
   234 => x"49d1c1f0",
   235 => x"c487edf5",
   236 => x"05987086",
   237 => x"c0c887cd",
   238 => x"4966cc1e",
   239 => x"c487f8fd",
   240 => x"ff4b7086",
   241 => x"78c248d0",
   242 => x"cbf54873",
   243 => x"5b5e0e87",
   244 => x"c00e5d5c",
   245 => x"f0ffc01e",
   246 => x"f449c9c1",
   247 => x"1ed287fe",
   248 => x"49d0e4c2",
   249 => x"c887d0fd",
   250 => x"c14cc086",
   251 => x"acb7d284",
   252 => x"c287f804",
   253 => x"bf97d0e4",
   254 => x"99c0c349",
   255 => x"05a9c0c1",
   256 => x"c287e7c0",
   257 => x"bf97d7e4",
   258 => x"c231d049",
   259 => x"bf97d8e4",
   260 => x"7232c84a",
   261 => x"d9e4c2b1",
   262 => x"b14abf97",
   263 => x"ffcf4c71",
   264 => x"c19cffff",
   265 => x"c134ca84",
   266 => x"e4c287e7",
   267 => x"49bf97d9",
   268 => x"99c631c1",
   269 => x"97dae4c2",
   270 => x"b7c74abf",
   271 => x"c2b1722a",
   272 => x"bf97d5e4",
   273 => x"9dcf4d4a",
   274 => x"97d6e4c2",
   275 => x"9ac34abf",
   276 => x"e4c232ca",
   277 => x"4bbf97d7",
   278 => x"b27333c2",
   279 => x"97d8e4c2",
   280 => x"c0c34bbf",
   281 => x"2bb7c69b",
   282 => x"81c2b273",
   283 => x"307148c1",
   284 => x"48c14970",
   285 => x"4d703075",
   286 => x"84c14c72",
   287 => x"c0c89471",
   288 => x"cc06adb7",
   289 => x"b734c187",
   290 => x"b7c0c82d",
   291 => x"f4ff01ad",
   292 => x"f1487487",
   293 => x"5e0e87fe",
   294 => x"0e5d5c5b",
   295 => x"ecc286f8",
   296 => x"78c048f6",
   297 => x"1eeee4c2",
   298 => x"defb49c0",
   299 => x"7086c487",
   300 => x"87c50598",
   301 => x"cec948c0",
   302 => x"c14dc087",
   303 => x"caf5c07e",
   304 => x"e5c249bf",
   305 => x"c8714ae4",
   306 => x"87deee4b",
   307 => x"c2059870",
   308 => x"c07ec087",
   309 => x"49bfc6f5",
   310 => x"4ac0e6c2",
   311 => x"ee4bc871",
   312 => x"987087c8",
   313 => x"c087c205",
   314 => x"c0026e7e",
   315 => x"ebc287fd",
   316 => x"c24dbff4",
   317 => x"bf9fecec",
   318 => x"d6c5487e",
   319 => x"c705a8ea",
   320 => x"f4ebc287",
   321 => x"87ce4dbf",
   322 => x"e9ca486e",
   323 => x"c502a8d5",
   324 => x"c748c087",
   325 => x"e4c287f1",
   326 => x"49751eee",
   327 => x"c487ecf9",
   328 => x"05987086",
   329 => x"48c087c5",
   330 => x"c087dcc7",
   331 => x"49bfc6f5",
   332 => x"4ac0e6c2",
   333 => x"ec4bc871",
   334 => x"987087f0",
   335 => x"c287c805",
   336 => x"c148f6ec",
   337 => x"c087da78",
   338 => x"49bfcaf5",
   339 => x"4ae4e5c2",
   340 => x"ec4bc871",
   341 => x"987087d4",
   342 => x"87c5c002",
   343 => x"e6c648c0",
   344 => x"ececc287",
   345 => x"c149bf97",
   346 => x"c005a9d5",
   347 => x"ecc287cd",
   348 => x"49bf97ed",
   349 => x"02a9eac2",
   350 => x"c087c5c0",
   351 => x"87c7c648",
   352 => x"97eee4c2",
   353 => x"c3487ebf",
   354 => x"c002a8e9",
   355 => x"486e87ce",
   356 => x"02a8ebc3",
   357 => x"c087c5c0",
   358 => x"87ebc548",
   359 => x"97f9e4c2",
   360 => x"059949bf",
   361 => x"c287ccc0",
   362 => x"bf97fae4",
   363 => x"02a9c249",
   364 => x"c087c5c0",
   365 => x"87cfc548",
   366 => x"97fbe4c2",
   367 => x"ecc248bf",
   368 => x"4c7058f2",
   369 => x"c288c148",
   370 => x"c258f6ec",
   371 => x"bf97fce4",
   372 => x"c2817549",
   373 => x"bf97fde4",
   374 => x"7232c84a",
   375 => x"f1c27ea1",
   376 => x"786e48c3",
   377 => x"97fee4c2",
   378 => x"a6c848bf",
   379 => x"f6ecc258",
   380 => x"d4c202bf",
   381 => x"c6f5c087",
   382 => x"e6c249bf",
   383 => x"c8714ac0",
   384 => x"87e6e94b",
   385 => x"c0029870",
   386 => x"48c087c5",
   387 => x"c287f8c3",
   388 => x"4cbfeeec",
   389 => x"5cd7f1c2",
   390 => x"97d3e5c2",
   391 => x"31c849bf",
   392 => x"97d2e5c2",
   393 => x"49a14abf",
   394 => x"97d4e5c2",
   395 => x"32d04abf",
   396 => x"c249a172",
   397 => x"bf97d5e5",
   398 => x"7232d84a",
   399 => x"66c449a1",
   400 => x"c3f1c291",
   401 => x"f1c281bf",
   402 => x"e5c259cb",
   403 => x"4abf97db",
   404 => x"e5c232c8",
   405 => x"4bbf97da",
   406 => x"e5c24aa2",
   407 => x"4bbf97dc",
   408 => x"a27333d0",
   409 => x"dde5c24a",
   410 => x"cf4bbf97",
   411 => x"7333d89b",
   412 => x"f1c24aa2",
   413 => x"f1c25acf",
   414 => x"c24abfcb",
   415 => x"c292748a",
   416 => x"7248cff1",
   417 => x"cac178a1",
   418 => x"c0e5c287",
   419 => x"c849bf97",
   420 => x"ffe4c231",
   421 => x"a14abf97",
   422 => x"feecc249",
   423 => x"faecc259",
   424 => x"31c549bf",
   425 => x"c981ffc7",
   426 => x"d7f1c229",
   427 => x"c5e5c259",
   428 => x"c84abf97",
   429 => x"c4e5c232",
   430 => x"a24bbf97",
   431 => x"9266c44a",
   432 => x"f1c2826e",
   433 => x"f1c25ad3",
   434 => x"78c048cb",
   435 => x"48c7f1c2",
   436 => x"c278a172",
   437 => x"c248d7f1",
   438 => x"78bfcbf1",
   439 => x"48dbf1c2",
   440 => x"bfcff1c2",
   441 => x"f6ecc278",
   442 => x"c9c002bf",
   443 => x"c4487487",
   444 => x"c07e7030",
   445 => x"f1c287c9",
   446 => x"c448bfd3",
   447 => x"c27e7030",
   448 => x"6e48faec",
   449 => x"f848c178",
   450 => x"264d268e",
   451 => x"264b264c",
   452 => x"5b5e0e4f",
   453 => x"710e5d5c",
   454 => x"f6ecc24a",
   455 => x"87cb02bf",
   456 => x"2bc74b72",
   457 => x"ffc14c72",
   458 => x"7287c99c",
   459 => x"722bc84b",
   460 => x"9cffc34c",
   461 => x"bfc3f1c2",
   462 => x"c2f5c083",
   463 => x"d902abbf",
   464 => x"c6f5c087",
   465 => x"eee4c25b",
   466 => x"f049731e",
   467 => x"86c487fd",
   468 => x"c5059870",
   469 => x"c048c087",
   470 => x"ecc287e6",
   471 => x"d202bff6",
   472 => x"c4497487",
   473 => x"eee4c291",
   474 => x"cf4d6981",
   475 => x"ffffffff",
   476 => x"7487cb9d",
   477 => x"c291c249",
   478 => x"9f81eee4",
   479 => x"48754d69",
   480 => x"0e87c6fe",
   481 => x"5d5c5b5e",
   482 => x"4d711e0e",
   483 => x"49c11ec0",
   484 => x"c487d7cf",
   485 => x"9c4c7086",
   486 => x"87c0c102",
   487 => x"4afeecc2",
   488 => x"eae24975",
   489 => x"02987087",
   490 => x"7487f1c0",
   491 => x"cb49754a",
   492 => x"87d0e34b",
   493 => x"c0029870",
   494 => x"1ec087e2",
   495 => x"c7029c74",
   496 => x"48a6c487",
   497 => x"87c578c0",
   498 => x"c148a6c4",
   499 => x"4966c478",
   500 => x"c487d7ce",
   501 => x"9c4c7086",
   502 => x"87c0ff05",
   503 => x"fc264874",
   504 => x"5e0e87e7",
   505 => x"0e5d5c5b",
   506 => x"9b4b711e",
   507 => x"c087c505",
   508 => x"87e5c148",
   509 => x"c04da3c8",
   510 => x"0266d47d",
   511 => x"66d487c7",
   512 => x"c505bf97",
   513 => x"c148c087",
   514 => x"66d487cf",
   515 => x"87f3fd49",
   516 => x"029c4c70",
   517 => x"dc87c0c1",
   518 => x"7d6949a4",
   519 => x"c449a4da",
   520 => x"699f4aa3",
   521 => x"f6ecc27a",
   522 => x"87d202bf",
   523 => x"9f49a4d4",
   524 => x"ffc04969",
   525 => x"487199ff",
   526 => x"7e7030d0",
   527 => x"7ec087c2",
   528 => x"6a48496e",
   529 => x"c07a7080",
   530 => x"49a3cc7b",
   531 => x"a3d0796a",
   532 => x"7479c049",
   533 => x"c087c248",
   534 => x"ecfa2648",
   535 => x"5b5e0e87",
   536 => x"710e5d5c",
   537 => x"c2f5c04c",
   538 => x"7478ff48",
   539 => x"cac1029c",
   540 => x"49a4c887",
   541 => x"c2c10269",
   542 => x"4a66d087",
   543 => x"d482496c",
   544 => x"66d05aa6",
   545 => x"ecc2b94d",
   546 => x"ff4abff2",
   547 => x"719972ba",
   548 => x"e4c00299",
   549 => x"4ba4c487",
   550 => x"f4f9496b",
   551 => x"c27b7087",
   552 => x"49bfeeec",
   553 => x"7c71816c",
   554 => x"ecc2b975",
   555 => x"ff4abff2",
   556 => x"719972ba",
   557 => x"dcff0599",
   558 => x"f97c7587",
   559 => x"731e87cb",
   560 => x"9b4b711e",
   561 => x"c887c702",
   562 => x"056949a3",
   563 => x"48c087c5",
   564 => x"c287ebc0",
   565 => x"4abfc7f1",
   566 => x"6949a3c4",
   567 => x"c289c249",
   568 => x"91bfeeec",
   569 => x"c24aa271",
   570 => x"49bff2ec",
   571 => x"a271996b",
   572 => x"1e66c84a",
   573 => x"d2ea4972",
   574 => x"7086c487",
   575 => x"ccf84849",
   576 => x"5b5e0e87",
   577 => x"1e0e5d5c",
   578 => x"66d44b71",
   579 => x"732cc94c",
   580 => x"cfc1029b",
   581 => x"49a3c887",
   582 => x"c7c10269",
   583 => x"4da3d087",
   584 => x"c27d66d4",
   585 => x"49bff2ec",
   586 => x"4a6bb9ff",
   587 => x"ac717e99",
   588 => x"c087cd03",
   589 => x"a3cc7d7b",
   590 => x"49a3c44a",
   591 => x"87c2796a",
   592 => x"9c748c72",
   593 => x"4987dd02",
   594 => x"fc49731e",
   595 => x"86c487cf",
   596 => x"c74966d4",
   597 => x"cb0299ff",
   598 => x"eee4c287",
   599 => x"fd49731e",
   600 => x"86c487dc",
   601 => x"87e1f626",
   602 => x"5c5b5e0e",
   603 => x"86f00e5d",
   604 => x"c059a6d0",
   605 => x"cc4b66e4",
   606 => x"87ca0266",
   607 => x"7080c848",
   608 => x"05bf6e7e",
   609 => x"48c087c5",
   610 => x"cc87ecc3",
   611 => x"84d04c66",
   612 => x"a6c44973",
   613 => x"c4786c48",
   614 => x"80c48166",
   615 => x"c878bf6e",
   616 => x"c606a966",
   617 => x"66c44987",
   618 => x"c04b7189",
   619 => x"c401abb7",
   620 => x"c2c34887",
   621 => x"4866c487",
   622 => x"7098ffc7",
   623 => x"c1026e7e",
   624 => x"c0c887c9",
   625 => x"71896e49",
   626 => x"eee4c24a",
   627 => x"73856e4d",
   628 => x"c106aab7",
   629 => x"49724a87",
   630 => x"8066c448",
   631 => x"8b727c70",
   632 => x"718ac149",
   633 => x"87d90299",
   634 => x"4866e0c0",
   635 => x"e0c05015",
   636 => x"80c14866",
   637 => x"58a6e4c0",
   638 => x"8ac14972",
   639 => x"e7059971",
   640 => x"d01ec187",
   641 => x"d4f94966",
   642 => x"c086c487",
   643 => x"c106abb7",
   644 => x"e0c087e3",
   645 => x"ffc74d66",
   646 => x"c006abb7",
   647 => x"1e7587e2",
   648 => x"fa4966d0",
   649 => x"c0c887d8",
   650 => x"c8486c85",
   651 => x"7c7080c0",
   652 => x"c18bc0c8",
   653 => x"4966d41e",
   654 => x"c887e2f8",
   655 => x"87eec086",
   656 => x"1eeee4c2",
   657 => x"f94966d0",
   658 => x"86c487f4",
   659 => x"4aeee4c2",
   660 => x"6c484973",
   661 => x"737c7080",
   662 => x"718bc149",
   663 => x"87ce0299",
   664 => x"c17d9712",
   665 => x"c1497385",
   666 => x"0599718b",
   667 => x"b7c087f2",
   668 => x"e1fe01ab",
   669 => x"f048c187",
   670 => x"87cdf28e",
   671 => x"5c5b5e0e",
   672 => x"4b710e5d",
   673 => x"87c7029b",
   674 => x"6d4da3c8",
   675 => x"ff87c505",
   676 => x"87fdc048",
   677 => x"6c4ca3d0",
   678 => x"99ffc749",
   679 => x"6c87d805",
   680 => x"c187c902",
   681 => x"f649731e",
   682 => x"86c487f3",
   683 => x"1eeee4c2",
   684 => x"c9f84973",
   685 => x"6c86c487",
   686 => x"04aa6d4a",
   687 => x"48ff87c4",
   688 => x"a2c187cf",
   689 => x"c749727c",
   690 => x"e4c299ff",
   691 => x"699781ee",
   692 => x"87f5f048",
   693 => x"711e731e",
   694 => x"c0029b4b",
   695 => x"f1c287e4",
   696 => x"4a735bdb",
   697 => x"ecc28ac2",
   698 => x"9249bfee",
   699 => x"bfc7f1c2",
   700 => x"c2807248",
   701 => x"7158dff1",
   702 => x"c230c448",
   703 => x"c058feec",
   704 => x"f1c287ed",
   705 => x"f1c248d7",
   706 => x"c278bfcb",
   707 => x"c248dbf1",
   708 => x"78bfcff1",
   709 => x"bff6ecc2",
   710 => x"c287c902",
   711 => x"49bfeeec",
   712 => x"87c731c4",
   713 => x"bfd3f1c2",
   714 => x"c231c449",
   715 => x"ef59feec",
   716 => x"5e0e87db",
   717 => x"710e5c5b",
   718 => x"724bc04a",
   719 => x"e1c0029a",
   720 => x"49a2da87",
   721 => x"c24b699f",
   722 => x"02bff6ec",
   723 => x"a2d487cf",
   724 => x"49699f49",
   725 => x"ffffc04c",
   726 => x"c234d09c",
   727 => x"744cc087",
   728 => x"4973b349",
   729 => x"ee87edfd",
   730 => x"5e0e87e1",
   731 => x"0e5d5c5b",
   732 => x"4a7186f4",
   733 => x"9a727ec0",
   734 => x"c287d802",
   735 => x"c048eae4",
   736 => x"e2e4c278",
   737 => x"dbf1c248",
   738 => x"e4c278bf",
   739 => x"f1c248e6",
   740 => x"c278bfd7",
   741 => x"c048cbed",
   742 => x"faecc250",
   743 => x"e4c249bf",
   744 => x"714abfea",
   745 => x"c0c403aa",
   746 => x"cf497287",
   747 => x"e1c00599",
   748 => x"eee4c287",
   749 => x"e2e4c21e",
   750 => x"e4c249bf",
   751 => x"a1c148e2",
   752 => x"dfff7178",
   753 => x"86c487c5",
   754 => x"48fef4c0",
   755 => x"78eee4c2",
   756 => x"f4c087cc",
   757 => x"c048bffe",
   758 => x"f5c080e0",
   759 => x"e4c258c2",
   760 => x"c148bfea",
   761 => x"eee4c280",
   762 => x"0d3e2758",
   763 => x"97bf0000",
   764 => x"029d4dbf",
   765 => x"c387e2c2",
   766 => x"c202ade5",
   767 => x"f4c087db",
   768 => x"cb4bbffe",
   769 => x"4c1149a3",
   770 => x"c105accf",
   771 => x"497587d2",
   772 => x"89c199df",
   773 => x"ecc291cd",
   774 => x"a3c181fe",
   775 => x"c351124a",
   776 => x"51124aa3",
   777 => x"124aa3c5",
   778 => x"4aa3c751",
   779 => x"a3c95112",
   780 => x"ce51124a",
   781 => x"51124aa3",
   782 => x"124aa3d0",
   783 => x"4aa3d251",
   784 => x"a3d45112",
   785 => x"d651124a",
   786 => x"51124aa3",
   787 => x"124aa3d8",
   788 => x"4aa3dc51",
   789 => x"a3de5112",
   790 => x"c151124a",
   791 => x"87f9c07e",
   792 => x"99c84974",
   793 => x"87eac005",
   794 => x"99d04974",
   795 => x"dc87d005",
   796 => x"cac00266",
   797 => x"dc497387",
   798 => x"98700f66",
   799 => x"6e87d302",
   800 => x"87c6c005",
   801 => x"48feecc2",
   802 => x"f4c050c0",
   803 => x"c248bffe",
   804 => x"edc287e7",
   805 => x"50c048cb",
   806 => x"faecc27e",
   807 => x"e4c249bf",
   808 => x"714abfea",
   809 => x"c0fc04aa",
   810 => x"dbf1c287",
   811 => x"c8c005bf",
   812 => x"f6ecc287",
   813 => x"fec102bf",
   814 => x"c2f5c087",
   815 => x"c278ff48",
   816 => x"49bfe6e4",
   817 => x"7087cae9",
   818 => x"eae4c249",
   819 => x"48a6c459",
   820 => x"bfe6e4c2",
   821 => x"f6ecc278",
   822 => x"d8c002bf",
   823 => x"4966c487",
   824 => x"ffffffcf",
   825 => x"02a999f8",
   826 => x"c087c5c0",
   827 => x"87e1c04d",
   828 => x"dcc04dc1",
   829 => x"4966c487",
   830 => x"99f8ffcf",
   831 => x"c8c002a9",
   832 => x"48a6c887",
   833 => x"c5c078c0",
   834 => x"48a6c887",
   835 => x"66c878c1",
   836 => x"059d754d",
   837 => x"c487e0c0",
   838 => x"89c24966",
   839 => x"bfeeecc2",
   840 => x"f1c2914a",
   841 => x"c24abfc7",
   842 => x"7248e2e4",
   843 => x"e4c278a1",
   844 => x"78c048ea",
   845 => x"c087e2f9",
   846 => x"e78ef448",
   847 => x"000087cb",
   848 => x"ffff0000",
   849 => x"0d4effff",
   850 => x"0d570000",
   851 => x"41460000",
   852 => x"20323354",
   853 => x"46002020",
   854 => x"36315441",
   855 => x"00202020",
   856 => x"e0f1c21e",
   857 => x"a8dd48bf",
   858 => x"c087c905",
   859 => x"7087d0ff",
   860 => x"87c84a49",
   861 => x"c348d4ff",
   862 => x"4a6878ff",
   863 => x"4f264872",
   864 => x"e0f1c21e",
   865 => x"a8dd48bf",
   866 => x"c087c605",
   867 => x"d987dcfe",
   868 => x"48d4ff87",
   869 => x"ff78ffc3",
   870 => x"e1c848d0",
   871 => x"48d4ff78",
   872 => x"f1c278d4",
   873 => x"d4ff48df",
   874 => x"4f2650bf",
   875 => x"48d0ff1e",
   876 => x"2678e0c0",
   877 => x"e7fe1e4f",
   878 => x"99497087",
   879 => x"c087c602",
   880 => x"f105a9fb",
   881 => x"26487187",
   882 => x"5b5e0e4f",
   883 => x"4b710e5c",
   884 => x"cbfe4cc0",
   885 => x"99497087",
   886 => x"87f9c002",
   887 => x"02a9ecc0",
   888 => x"c087f2c0",
   889 => x"c002a9fb",
   890 => x"66cc87eb",
   891 => x"c703acb7",
   892 => x"0266d087",
   893 => x"537187c2",
   894 => x"c2029971",
   895 => x"fd84c187",
   896 => x"497087de",
   897 => x"87cd0299",
   898 => x"02a9ecc0",
   899 => x"fbc087c7",
   900 => x"d5ff05a9",
   901 => x"0266d087",
   902 => x"97c087c3",
   903 => x"a9ecc07b",
   904 => x"7487c405",
   905 => x"7487c54a",
   906 => x"8a0ac04a",
   907 => x"87c24872",
   908 => x"4c264d26",
   909 => x"4f264b26",
   910 => x"87e4fc1e",
   911 => x"f0c04970",
   912 => x"ca04a9b7",
   913 => x"b7f9c087",
   914 => x"87c301a9",
   915 => x"c189f0c0",
   916 => x"04a9b7c1",
   917 => x"dac187ca",
   918 => x"c301a9b7",
   919 => x"89f7c087",
   920 => x"4f264871",
   921 => x"5c5b5e0e",
   922 => x"ff4a710e",
   923 => x"49724cd4",
   924 => x"7087eac0",
   925 => x"c2029b4b",
   926 => x"ff8bc187",
   927 => x"c5c848d0",
   928 => x"7cd5c178",
   929 => x"31c64973",
   930 => x"97f4e2c2",
   931 => x"71484abf",
   932 => x"ff7c70b0",
   933 => x"78c448d0",
   934 => x"d5fe4873",
   935 => x"5b5e0e87",
   936 => x"f40e5d5c",
   937 => x"c44c7186",
   938 => x"78c048a6",
   939 => x"6e7ea4c8",
   940 => x"c149bf97",
   941 => x"dd05a9c1",
   942 => x"49a4c987",
   943 => x"c1496997",
   944 => x"d105a9d2",
   945 => x"49a4ca87",
   946 => x"c1496997",
   947 => x"c505a9c3",
   948 => x"c248df87",
   949 => x"e7fa87e1",
   950 => x"c04bc087",
   951 => x"bf97fcfd",
   952 => x"04a9c049",
   953 => x"ccfb87cf",
   954 => x"c083c187",
   955 => x"bf97fcfd",
   956 => x"f106ab49",
   957 => x"fcfdc087",
   958 => x"cf02bf97",
   959 => x"87e0f987",
   960 => x"02994970",
   961 => x"ecc087c6",
   962 => x"87f105a9",
   963 => x"cff94bc0",
   964 => x"f94d7087",
   965 => x"a6cc87ca",
   966 => x"87c4f958",
   967 => x"83c14a70",
   968 => x"49bf976e",
   969 => x"87c702ad",
   970 => x"05adffc0",
   971 => x"c987eac0",
   972 => x"699749a4",
   973 => x"a966c849",
   974 => x"4887c702",
   975 => x"05a8ffc0",
   976 => x"a4ca87d7",
   977 => x"49699749",
   978 => x"87c602aa",
   979 => x"05aaffc0",
   980 => x"a6c487c7",
   981 => x"d378c148",
   982 => x"adecc087",
   983 => x"c087c602",
   984 => x"c705adfb",
   985 => x"c44bc087",
   986 => x"78c148a6",
   987 => x"fe0266c4",
   988 => x"f7f887dc",
   989 => x"f4487387",
   990 => x"87f4fa8e",
   991 => x"5b5e0e00",
   992 => x"1e0e5d5c",
   993 => x"4cc04b71",
   994 => x"c004ab4d",
   995 => x"fac087e8",
   996 => x"9d751edd",
   997 => x"c087c402",
   998 => x"c187c24a",
   999 => x"ef49724a",
  1000 => x"86c487c8",
  1001 => x"84c17e70",
  1002 => x"87c2056e",
  1003 => x"85c14c73",
  1004 => x"ff06ac73",
  1005 => x"486e87d8",
  1006 => x"264d2626",
  1007 => x"264b264c",
  1008 => x"5b5e0e4f",
  1009 => x"1e0e5d5c",
  1010 => x"de494c71",
  1011 => x"f9f1c291",
  1012 => x"9785714d",
  1013 => x"ddc1026d",
  1014 => x"e4f1c287",
  1015 => x"82744abf",
  1016 => x"d8fe4972",
  1017 => x"6e7e7087",
  1018 => x"87f3c002",
  1019 => x"4becf1c2",
  1020 => x"49cb4a6e",
  1021 => x"87f0c2ff",
  1022 => x"93cb4b74",
  1023 => x"83d0e2c1",
  1024 => x"c0c183c4",
  1025 => x"49747bfa",
  1026 => x"87fecdc1",
  1027 => x"f1c27b75",
  1028 => x"49bf97f8",
  1029 => x"ecf1c21e",
  1030 => x"c8e2c149",
  1031 => x"7486c487",
  1032 => x"e5cdc149",
  1033 => x"c149c087",
  1034 => x"c287c4cf",
  1035 => x"c048e0f1",
  1036 => x"dd49c178",
  1037 => x"fd2687cf",
  1038 => x"6f4c87ff",
  1039 => x"6e696461",
  1040 => x"2e2e2e67",
  1041 => x"5b5e0e00",
  1042 => x"4b710e5c",
  1043 => x"e4f1c24a",
  1044 => x"497282bf",
  1045 => x"7087e6fc",
  1046 => x"c4029c4c",
  1047 => x"d1eb4987",
  1048 => x"e4f1c287",
  1049 => x"c178c048",
  1050 => x"87d9dc49",
  1051 => x"0e87ccfd",
  1052 => x"5d5c5b5e",
  1053 => x"c286f40e",
  1054 => x"c04deee4",
  1055 => x"48a6c44c",
  1056 => x"f1c278c0",
  1057 => x"c049bfe4",
  1058 => x"c1c106a9",
  1059 => x"eee4c287",
  1060 => x"c0029848",
  1061 => x"fac087f8",
  1062 => x"66c81edd",
  1063 => x"c487c702",
  1064 => x"78c048a6",
  1065 => x"a6c487c5",
  1066 => x"c478c148",
  1067 => x"f9ea4966",
  1068 => x"7086c487",
  1069 => x"c484c14d",
  1070 => x"80c14866",
  1071 => x"c258a6c8",
  1072 => x"49bfe4f1",
  1073 => x"87c603ac",
  1074 => x"ff059d75",
  1075 => x"4cc087c8",
  1076 => x"c3029d75",
  1077 => x"fac087e0",
  1078 => x"66c81edd",
  1079 => x"cc87c702",
  1080 => x"78c048a6",
  1081 => x"a6cc87c5",
  1082 => x"cc78c148",
  1083 => x"f9e94966",
  1084 => x"7086c487",
  1085 => x"c2026e7e",
  1086 => x"496e87e9",
  1087 => x"699781cb",
  1088 => x"0299d049",
  1089 => x"c187d6c1",
  1090 => x"744ac5c1",
  1091 => x"c191cb49",
  1092 => x"7281d0e2",
  1093 => x"c381c879",
  1094 => x"497451ff",
  1095 => x"f1c291de",
  1096 => x"85714df9",
  1097 => x"7d97c1c2",
  1098 => x"c049a5c1",
  1099 => x"ecc251e0",
  1100 => x"02bf97fe",
  1101 => x"84c187d2",
  1102 => x"c24ba5c2",
  1103 => x"db4afeec",
  1104 => x"e3fdfe49",
  1105 => x"87dbc187",
  1106 => x"c049a5cd",
  1107 => x"c284c151",
  1108 => x"4a6e4ba5",
  1109 => x"fdfe49cb",
  1110 => x"c6c187ce",
  1111 => x"c1ffc087",
  1112 => x"cb49744a",
  1113 => x"d0e2c191",
  1114 => x"c2797281",
  1115 => x"bf97feec",
  1116 => x"7487d802",
  1117 => x"c191de49",
  1118 => x"f9f1c284",
  1119 => x"c283714b",
  1120 => x"dd4afeec",
  1121 => x"dffcfe49",
  1122 => x"7487d887",
  1123 => x"c293de4b",
  1124 => x"cb83f9f1",
  1125 => x"51c049a3",
  1126 => x"6e7384c1",
  1127 => x"fe49cb4a",
  1128 => x"c487c5fc",
  1129 => x"80c14866",
  1130 => x"c758a6c8",
  1131 => x"c5c003ac",
  1132 => x"fc056e87",
  1133 => x"487487e0",
  1134 => x"fcf78ef4",
  1135 => x"1e731e87",
  1136 => x"cb494b71",
  1137 => x"d0e2c191",
  1138 => x"4aa1c881",
  1139 => x"48f4e2c2",
  1140 => x"a1c95012",
  1141 => x"fcfdc04a",
  1142 => x"ca501248",
  1143 => x"f8f1c281",
  1144 => x"c2501148",
  1145 => x"bf97f8f1",
  1146 => x"49c01e49",
  1147 => x"87f5dac1",
  1148 => x"48e0f1c2",
  1149 => x"49c178de",
  1150 => x"2687cad6",
  1151 => x"1e87fef6",
  1152 => x"cb494a71",
  1153 => x"d0e2c191",
  1154 => x"1181c881",
  1155 => x"e4f1c248",
  1156 => x"e4f1c258",
  1157 => x"c178c048",
  1158 => x"87e9d549",
  1159 => x"c01e4f26",
  1160 => x"cac7c149",
  1161 => x"1e4f2687",
  1162 => x"d2029971",
  1163 => x"e5e3c187",
  1164 => x"f750c048",
  1165 => x"ffc7c180",
  1166 => x"c9e2c140",
  1167 => x"c187ce78",
  1168 => x"c148e1e3",
  1169 => x"fc78c2e2",
  1170 => x"dec8c180",
  1171 => x"0e4f2678",
  1172 => x"0e5c5b5e",
  1173 => x"cb4a4c71",
  1174 => x"d0e2c192",
  1175 => x"49a2c882",
  1176 => x"974ba2c9",
  1177 => x"971e4b6b",
  1178 => x"ca1e4969",
  1179 => x"c0491282",
  1180 => x"c087ebe7",
  1181 => x"87cdd449",
  1182 => x"c4c14974",
  1183 => x"8ef887cc",
  1184 => x"1e87f8f4",
  1185 => x"4b711e73",
  1186 => x"87c3ff49",
  1187 => x"fefe4973",
  1188 => x"87e9f487",
  1189 => x"711e731e",
  1190 => x"4aa3c64b",
  1191 => x"c187db02",
  1192 => x"87d6028a",
  1193 => x"dac1028a",
  1194 => x"c0028a87",
  1195 => x"028a87fc",
  1196 => x"8a87e1c0",
  1197 => x"c187cb02",
  1198 => x"49c787db",
  1199 => x"c187c0fd",
  1200 => x"f1c287de",
  1201 => x"c102bfe4",
  1202 => x"c14887cb",
  1203 => x"e8f1c288",
  1204 => x"87c1c158",
  1205 => x"bfe8f1c2",
  1206 => x"87f9c002",
  1207 => x"bfe4f1c2",
  1208 => x"c280c148",
  1209 => x"c058e8f1",
  1210 => x"f1c287eb",
  1211 => x"c649bfe4",
  1212 => x"e8f1c289",
  1213 => x"a9b7c059",
  1214 => x"c287da03",
  1215 => x"c048e4f1",
  1216 => x"c287d278",
  1217 => x"02bfe8f1",
  1218 => x"f1c287cb",
  1219 => x"c648bfe4",
  1220 => x"e8f1c280",
  1221 => x"d149c058",
  1222 => x"497387eb",
  1223 => x"87eac1c1",
  1224 => x"1e87daf2",
  1225 => x"4b711e73",
  1226 => x"48e0f1c2",
  1227 => x"49c078dd",
  1228 => x"7387d2d1",
  1229 => x"d1c1c149",
  1230 => x"87c1f287",
  1231 => x"5c5b5e0e",
  1232 => x"cc4c710e",
  1233 => x"4b741e66",
  1234 => x"e2c193cb",
  1235 => x"a3c483d0",
  1236 => x"fe496a4a",
  1237 => x"c187e1f5",
  1238 => x"c87bfdc6",
  1239 => x"66d449a3",
  1240 => x"49a3c951",
  1241 => x"ca5166d8",
  1242 => x"66dc49a3",
  1243 => x"caf12651",
  1244 => x"5b5e0e87",
  1245 => x"ff0e5d5c",
  1246 => x"a6dc86cc",
  1247 => x"48a6c859",
  1248 => x"80c478c0",
  1249 => x"7866c8c1",
  1250 => x"78c180c4",
  1251 => x"78c180c4",
  1252 => x"48e8f1c2",
  1253 => x"f1c278c1",
  1254 => x"de48bfe0",
  1255 => x"87cb05a8",
  1256 => x"7087ccf3",
  1257 => x"59a6cc49",
  1258 => x"e787d6ce",
  1259 => x"c4e887d2",
  1260 => x"87ece687",
  1261 => x"fbc04c70",
  1262 => x"d8c102ac",
  1263 => x"0566d887",
  1264 => x"c087cac1",
  1265 => x"1ec11e1e",
  1266 => x"1ec3e4c1",
  1267 => x"ebfd49c0",
  1268 => x"c086d087",
  1269 => x"d902acfb",
  1270 => x"66c4c187",
  1271 => x"6a82c44a",
  1272 => x"7481c749",
  1273 => x"d81ec151",
  1274 => x"c8496a1e",
  1275 => x"87d9e781",
  1276 => x"c8c186c8",
  1277 => x"a8c04866",
  1278 => x"c887c701",
  1279 => x"78c148a6",
  1280 => x"c8c187ce",
  1281 => x"88c14866",
  1282 => x"c358a6d0",
  1283 => x"87e5e687",
  1284 => x"c248a6d0",
  1285 => x"029c7478",
  1286 => x"c887e2cc",
  1287 => x"ccc14866",
  1288 => x"cc03a866",
  1289 => x"a6dc87d7",
  1290 => x"e478c048",
  1291 => x"4c7087f2",
  1292 => x"dd4866d8",
  1293 => x"87c605a8",
  1294 => x"d848a6dc",
  1295 => x"d0c17866",
  1296 => x"e8c005ac",
  1297 => x"87d8e487",
  1298 => x"7087d5e4",
  1299 => x"acecc04c",
  1300 => x"e587c505",
  1301 => x"4c7087df",
  1302 => x"05acd0c1",
  1303 => x"66d487c8",
  1304 => x"d880c148",
  1305 => x"d0c158a6",
  1306 => x"d8ff02ac",
  1307 => x"a6e0c087",
  1308 => x"7866d848",
  1309 => x"c04866dc",
  1310 => x"05a866e0",
  1311 => x"c487d0ca",
  1312 => x"f0c048a6",
  1313 => x"80e0c078",
  1314 => x"c47866d0",
  1315 => x"c478c080",
  1316 => x"7478c080",
  1317 => x"8dfbc04d",
  1318 => x"87ccc902",
  1319 => x"db028dc9",
  1320 => x"028dc287",
  1321 => x"c987cdc1",
  1322 => x"d1c4028d",
  1323 => x"028dc487",
  1324 => x"c187cec1",
  1325 => x"c5c4028d",
  1326 => x"87e6c887",
  1327 => x"cb4966c8",
  1328 => x"66c4c191",
  1329 => x"4aa1c481",
  1330 => x"1e717e6a",
  1331 => x"48f8ddc1",
  1332 => x"cc4966c4",
  1333 => x"41204aa1",
  1334 => x"ff05aa71",
  1335 => x"511087f8",
  1336 => x"ccc14926",
  1337 => x"cce379e3",
  1338 => x"c04c7087",
  1339 => x"c148a6ec",
  1340 => x"87f4c778",
  1341 => x"c048a6c4",
  1342 => x"4866d078",
  1343 => x"a6d480c1",
  1344 => x"87dce158",
  1345 => x"ecc04c70",
  1346 => x"87d402ac",
  1347 => x"c00266c4",
  1348 => x"a6c887c5",
  1349 => x"7487c95c",
  1350 => x"88f0c048",
  1351 => x"58a6e8c0",
  1352 => x"02acecc0",
  1353 => x"f7e087cc",
  1354 => x"c04c7087",
  1355 => x"ff05acec",
  1356 => x"66c487f4",
  1357 => x"4966d81e",
  1358 => x"66ecc01e",
  1359 => x"c3e4c11e",
  1360 => x"4966d81e",
  1361 => x"c087f5f7",
  1362 => x"c01eca1e",
  1363 => x"cb4966e0",
  1364 => x"66dcc191",
  1365 => x"48a6d881",
  1366 => x"d878a1c4",
  1367 => x"e149bf66",
  1368 => x"86d887e7",
  1369 => x"06a8b7c0",
  1370 => x"c187cac1",
  1371 => x"c81ede1e",
  1372 => x"e149bf66",
  1373 => x"86c887d3",
  1374 => x"c0484970",
  1375 => x"e8c08808",
  1376 => x"b7c058a6",
  1377 => x"ecc006a8",
  1378 => x"66e4c087",
  1379 => x"a8b7dd48",
  1380 => x"87e1c003",
  1381 => x"c049bf6e",
  1382 => x"c08166e4",
  1383 => x"e4c051e0",
  1384 => x"81c14966",
  1385 => x"c281bf6e",
  1386 => x"e4c051c1",
  1387 => x"81c24966",
  1388 => x"c081bf6e",
  1389 => x"a6ecc051",
  1390 => x"c478c148",
  1391 => x"f7e187ea",
  1392 => x"a6e8c087",
  1393 => x"87f0e158",
  1394 => x"58a6f0c0",
  1395 => x"05a8ecc0",
  1396 => x"a687c9c0",
  1397 => x"66e4c048",
  1398 => x"87c4c078",
  1399 => x"87c0deff",
  1400 => x"cb4966c8",
  1401 => x"66c4c191",
  1402 => x"c8807148",
  1403 => x"66c458a6",
  1404 => x"c482c84a",
  1405 => x"81ca4966",
  1406 => x"5166e4c0",
  1407 => x"4966ecc0",
  1408 => x"e4c081c1",
  1409 => x"48c18966",
  1410 => x"49703071",
  1411 => x"977189c1",
  1412 => x"d5f5c27a",
  1413 => x"e4c049bf",
  1414 => x"6a972966",
  1415 => x"9871484a",
  1416 => x"58a6f4c0",
  1417 => x"c44966c4",
  1418 => x"c07e6981",
  1419 => x"dc4866e0",
  1420 => x"c002a866",
  1421 => x"a6dc87c8",
  1422 => x"c078c048",
  1423 => x"a6dc87c5",
  1424 => x"dc78c148",
  1425 => x"e0c01e66",
  1426 => x"4966c81e",
  1427 => x"87f9ddff",
  1428 => x"4c7086c8",
  1429 => x"06acb7c0",
  1430 => x"6e87d6c1",
  1431 => x"70807448",
  1432 => x"49e0c07e",
  1433 => x"4b6e8974",
  1434 => x"4af5ddc1",
  1435 => x"f7e8fe71",
  1436 => x"c2486e87",
  1437 => x"c07e7080",
  1438 => x"c14866e8",
  1439 => x"a6ecc080",
  1440 => x"66f0c058",
  1441 => x"7081c149",
  1442 => x"c5c002a9",
  1443 => x"c04dc087",
  1444 => x"4dc187c2",
  1445 => x"a4c21e75",
  1446 => x"48e0c049",
  1447 => x"49708871",
  1448 => x"4966c81e",
  1449 => x"87e1dcff",
  1450 => x"b7c086c8",
  1451 => x"c6ff01a8",
  1452 => x"66e8c087",
  1453 => x"87d3c002",
  1454 => x"c94966c4",
  1455 => x"66e8c081",
  1456 => x"4866c451",
  1457 => x"78cfc9c1",
  1458 => x"c487cec0",
  1459 => x"81c94966",
  1460 => x"66c451c2",
  1461 => x"c3cac148",
  1462 => x"a6ecc078",
  1463 => x"c078c148",
  1464 => x"dbff87c6",
  1465 => x"4c7087cf",
  1466 => x"0266ecc0",
  1467 => x"c887f5c0",
  1468 => x"66cc4866",
  1469 => x"cbc004a8",
  1470 => x"4866c887",
  1471 => x"a6cc80c1",
  1472 => x"87e0c058",
  1473 => x"c14866cc",
  1474 => x"58a6d088",
  1475 => x"c187d5c0",
  1476 => x"c005acc6",
  1477 => x"66d087c8",
  1478 => x"d480c148",
  1479 => x"daff58a6",
  1480 => x"4c7087d3",
  1481 => x"c14866d4",
  1482 => x"58a6d880",
  1483 => x"c0029c74",
  1484 => x"66c887cb",
  1485 => x"66ccc148",
  1486 => x"e9f304a8",
  1487 => x"ebd9ff87",
  1488 => x"4866c887",
  1489 => x"c003a8c7",
  1490 => x"f1c287e5",
  1491 => x"78c048e8",
  1492 => x"cb4966c8",
  1493 => x"66c4c191",
  1494 => x"4aa1c481",
  1495 => x"52c04a6a",
  1496 => x"4866c879",
  1497 => x"a6cc80c1",
  1498 => x"04a8c758",
  1499 => x"ff87dbff",
  1500 => x"c4e18ecc",
  1501 => x"00203a87",
  1502 => x"20504944",
  1503 => x"74697753",
  1504 => x"73656863",
  1505 => x"1e731e00",
  1506 => x"029b4b71",
  1507 => x"f1c287c6",
  1508 => x"78c048e4",
  1509 => x"f1c21ec7",
  1510 => x"1e49bfe4",
  1511 => x"1ed0e2c1",
  1512 => x"bfe0f1c2",
  1513 => x"87c9ef49",
  1514 => x"f1c286cc",
  1515 => x"e949bfe0",
  1516 => x"9b7387f5",
  1517 => x"c187c802",
  1518 => x"c049d0e2",
  1519 => x"ff87ddf0",
  1520 => x"1e87fadf",
  1521 => x"4bc01e73",
  1522 => x"48f4e2c2",
  1523 => x"e3c150c0",
  1524 => x"c049bff3",
  1525 => x"7087e5fe",
  1526 => x"87c40598",
  1527 => x"4be6dfc1",
  1528 => x"dfff4873",
  1529 => x"4f5287d7",
  1530 => x"6f6c204d",
  1531 => x"6e696461",
  1532 => x"61662067",
  1533 => x"64656c69",
  1534 => x"e5c71e00",
  1535 => x"fe49c187",
  1536 => x"eafe87c3",
  1537 => x"987087ec",
  1538 => x"fe87cd02",
  1539 => x"7087c7f2",
  1540 => x"87c40298",
  1541 => x"87c24ac1",
  1542 => x"9a724ac0",
  1543 => x"c087ce05",
  1544 => x"cde1c11e",
  1545 => x"d1fbc049",
  1546 => x"fe86c487",
  1547 => x"edc2c187",
  1548 => x"c11ec087",
  1549 => x"c049d8e1",
  1550 => x"c087fffa",
  1551 => x"87c3fe1e",
  1552 => x"fac04970",
  1553 => x"d8c387f4",
  1554 => x"268ef887",
  1555 => x"2044534f",
  1556 => x"6c696166",
  1557 => x"002e6465",
  1558 => x"746f6f42",
  1559 => x"2e676e69",
  1560 => x"1e002e2e",
  1561 => x"87d5f2c0",
  1562 => x"4f2687fa",
  1563 => x"e4f1c21e",
  1564 => x"c278c048",
  1565 => x"c048e0f1",
  1566 => x"87fdfd78",
  1567 => x"48c087e5",
  1568 => x"20804f26",
  1569 => x"74697845",
  1570 => x"42208000",
  1571 => x"006b6361",
  1572 => x"000011ff",
  1573 => x"00002c79",
  1574 => x"ff000000",
  1575 => x"97000011",
  1576 => x"0000002c",
  1577 => x"11ff0000",
  1578 => x"2cb50000",
  1579 => x"00000000",
  1580 => x"0011ff00",
  1581 => x"002cd300",
  1582 => x"00000000",
  1583 => x"000011ff",
  1584 => x"00002cf1",
  1585 => x"ff000000",
  1586 => x"0f000011",
  1587 => x"0000002d",
  1588 => x"11ff0000",
  1589 => x"2d2d0000",
  1590 => x"00000000",
  1591 => x"0011ff00",
  1592 => x"00000000",
  1593 => x"00000000",
  1594 => x"00001294",
  1595 => x"00000000",
  1596 => x"f7000000",
  1597 => x"4d000018",
  1598 => x"20554e45",
  1599 => x"52202020",
  1600 => x"4c004d4f",
  1601 => x"2064616f",
  1602 => x"1e002e2a",
  1603 => x"c048f0fe",
  1604 => x"7909cd78",
  1605 => x"1e4f2609",
  1606 => x"bff0fe1e",
  1607 => x"2626487e",
  1608 => x"f0fe1e4f",
  1609 => x"2678c148",
  1610 => x"f0fe1e4f",
  1611 => x"2678c048",
  1612 => x"4a711e4f",
  1613 => x"265252c0",
  1614 => x"5b5e0e4f",
  1615 => x"f40e5d5c",
  1616 => x"974d7186",
  1617 => x"a5c17e6d",
  1618 => x"486c974c",
  1619 => x"6e58a6c8",
  1620 => x"a866c448",
  1621 => x"ff87c505",
  1622 => x"87e6c048",
  1623 => x"c287caff",
  1624 => x"6c9749a5",
  1625 => x"4ba3714b",
  1626 => x"974b6b97",
  1627 => x"486e7e6c",
  1628 => x"a6c880c1",
  1629 => x"cc98c758",
  1630 => x"977058a6",
  1631 => x"87e1fe7c",
  1632 => x"8ef44873",
  1633 => x"4c264d26",
  1634 => x"4f264b26",
  1635 => x"5c5b5e0e",
  1636 => x"7186f40e",
  1637 => x"4a66d84c",
  1638 => x"c29affc3",
  1639 => x"6c974ba4",
  1640 => x"49a17349",
  1641 => x"6c975172",
  1642 => x"c1486e7e",
  1643 => x"58a6c880",
  1644 => x"a6cc98c7",
  1645 => x"f4547058",
  1646 => x"87caff8e",
  1647 => x"e8fd1e1e",
  1648 => x"4abfe087",
  1649 => x"c0e0c049",
  1650 => x"87cb0299",
  1651 => x"f5c21e72",
  1652 => x"f7fe49cb",
  1653 => x"fc86c487",
  1654 => x"7e7087fd",
  1655 => x"2687c2fd",
  1656 => x"c21e4f26",
  1657 => x"fd49cbf5",
  1658 => x"e6c187c7",
  1659 => x"dafc49fc",
  1660 => x"87d9c587",
  1661 => x"5e0e4f26",
  1662 => x"0e5d5c5b",
  1663 => x"bfdef6c2",
  1664 => x"cae9c14a",
  1665 => x"724c49bf",
  1666 => x"fc4d71bc",
  1667 => x"4bc087db",
  1668 => x"99d04974",
  1669 => x"7587d502",
  1670 => x"7199d049",
  1671 => x"c11ec01e",
  1672 => x"734adcef",
  1673 => x"c0491282",
  1674 => x"86c887e4",
  1675 => x"832d2cc1",
  1676 => x"ff04abc8",
  1677 => x"e8fb87da",
  1678 => x"cae9c187",
  1679 => x"def6c248",
  1680 => x"4d2678bf",
  1681 => x"4b264c26",
  1682 => x"00004f26",
  1683 => x"ff1e0000",
  1684 => x"e1c848d0",
  1685 => x"48d4ff78",
  1686 => x"66c478c5",
  1687 => x"c387c302",
  1688 => x"66c878e0",
  1689 => x"ff87c602",
  1690 => x"f0c348d4",
  1691 => x"48d4ff78",
  1692 => x"d0ff7871",
  1693 => x"78e1c848",
  1694 => x"2678e0c0",
  1695 => x"5b5e0e4f",
  1696 => x"4c710e5c",
  1697 => x"49cbf5c2",
  1698 => x"7087eefa",
  1699 => x"aab7c04a",
  1700 => x"87e3c204",
  1701 => x"05aae0c3",
  1702 => x"edc187c9",
  1703 => x"78c148c0",
  1704 => x"c387d4c2",
  1705 => x"c905aaf0",
  1706 => x"fcecc187",
  1707 => x"c178c148",
  1708 => x"edc187f5",
  1709 => x"c702bfc0",
  1710 => x"c24b7287",
  1711 => x"87c2b3c0",
  1712 => x"9c744b72",
  1713 => x"c187d105",
  1714 => x"1ebffcec",
  1715 => x"bfc0edc1",
  1716 => x"fd49721e",
  1717 => x"86c887f8",
  1718 => x"bffcecc1",
  1719 => x"87e0c002",
  1720 => x"b7c44973",
  1721 => x"eec19129",
  1722 => x"4a7381dc",
  1723 => x"92c29acf",
  1724 => x"307248c1",
  1725 => x"baff4a70",
  1726 => x"98694872",
  1727 => x"87db7970",
  1728 => x"b7c44973",
  1729 => x"eec19129",
  1730 => x"4a7381dc",
  1731 => x"92c29acf",
  1732 => x"307248c3",
  1733 => x"69484a70",
  1734 => x"c17970b0",
  1735 => x"c048c0ed",
  1736 => x"fcecc178",
  1737 => x"c278c048",
  1738 => x"f849cbf5",
  1739 => x"4a7087cb",
  1740 => x"03aab7c0",
  1741 => x"c087ddfd",
  1742 => x"87c8fc48",
  1743 => x"00000000",
  1744 => x"00000000",
  1745 => x"494a711e",
  1746 => x"2687f2fc",
  1747 => x"4ac01e4f",
  1748 => x"91c44972",
  1749 => x"81dceec1",
  1750 => x"82c179c0",
  1751 => x"04aab7d0",
  1752 => x"4f2687ee",
  1753 => x"5c5b5e0e",
  1754 => x"4d710e5d",
  1755 => x"7587faf6",
  1756 => x"2ab7c44a",
  1757 => x"dceec192",
  1758 => x"cf4c7582",
  1759 => x"6a94c29c",
  1760 => x"2b744b49",
  1761 => x"48c29bc3",
  1762 => x"4c703074",
  1763 => x"4874bcff",
  1764 => x"7a709871",
  1765 => x"7387caf6",
  1766 => x"87e6fa48",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"25261e16",
  1784 => x"3e3d362e",
  1785 => x"48d0ff1e",
  1786 => x"7178e1c8",
  1787 => x"08d4ff48",
  1788 => x"4866c478",
  1789 => x"7808d4ff",
  1790 => x"711e4f26",
  1791 => x"4966c44a",
  1792 => x"ff49721e",
  1793 => x"d0ff87de",
  1794 => x"78e0c048",
  1795 => x"1e4f2626",
  1796 => x"66c44a71",
  1797 => x"a2e0c11e",
  1798 => x"87c8ff49",
  1799 => x"c84966c8",
  1800 => x"d4ff29b7",
  1801 => x"ff787148",
  1802 => x"e0c048d0",
  1803 => x"4f262678",
  1804 => x"4ad4ff1e",
  1805 => x"ff7affc3",
  1806 => x"e1c848d0",
  1807 => x"c27ade78",
  1808 => x"7abfd5f5",
  1809 => x"28c84849",
  1810 => x"48717a70",
  1811 => x"7a7028d0",
  1812 => x"28d84871",
  1813 => x"d0ff7a70",
  1814 => x"78e0c048",
  1815 => x"5e0e4f26",
  1816 => x"0e5d5c5b",
  1817 => x"f5c24c71",
  1818 => x"4b4dbfd5",
  1819 => x"66d02b74",
  1820 => x"d483c19b",
  1821 => x"c204ab66",
  1822 => x"744bc087",
  1823 => x"4966d04a",
  1824 => x"b9ff3172",
  1825 => x"48739975",
  1826 => x"4a703072",
  1827 => x"c2b07148",
  1828 => x"fe58d9f5",
  1829 => x"4d2687da",
  1830 => x"4b264c26",
  1831 => x"5e0e4f26",
  1832 => x"0e5d5c5b",
  1833 => x"c24c711e",
  1834 => x"c04bd9f5",
  1835 => x"49f4c04a",
  1836 => x"87d1d0fe",
  1837 => x"f5c21e74",
  1838 => x"ecfe49d9",
  1839 => x"86c487e4",
  1840 => x"c0029870",
  1841 => x"1ec487ea",
  1842 => x"c21e4da6",
  1843 => x"fe49d9f5",
  1844 => x"c887d5f2",
  1845 => x"02987086",
  1846 => x"4a7587d6",
  1847 => x"49e6f4c1",
  1848 => x"cefe4bc4",
  1849 => x"987087c4",
  1850 => x"c087ca02",
  1851 => x"87edc048",
  1852 => x"e8c048c0",
  1853 => x"87f3c087",
  1854 => x"7087c4c1",
  1855 => x"87c80298",
  1856 => x"7087fcc0",
  1857 => x"87f80598",
  1858 => x"bff9f5c2",
  1859 => x"c287cc02",
  1860 => x"c248d5f5",
  1861 => x"78bff9f5",
  1862 => x"c187d5fc",
  1863 => x"4d262648",
  1864 => x"4b264c26",
  1865 => x"415b4f26",
  1866 => x"1e004352",
  1867 => x"f5c21ec0",
  1868 => x"effe49d9",
  1869 => x"f5c287cb",
  1870 => x"78c048f1",
  1871 => x"0e4f2626",
  1872 => x"5d5c5b5e",
  1873 => x"c486f40e",
  1874 => x"78c048a6",
  1875 => x"bff1f5c2",
  1876 => x"a8b7c348",
  1877 => x"c287d103",
  1878 => x"48bff1f5",
  1879 => x"f5c280c1",
  1880 => x"fbc058f5",
  1881 => x"87e2c648",
  1882 => x"49d9f5c2",
  1883 => x"87ccf4fe",
  1884 => x"f5c24c70",
  1885 => x"c34abff1",
  1886 => x"87d8028a",
  1887 => x"c5028ac1",
  1888 => x"028a87cb",
  1889 => x"8a87f6c2",
  1890 => x"87cdc102",
  1891 => x"e2c3028a",
  1892 => x"87e1c587",
  1893 => x"4a754dc0",
  1894 => x"fcc192c4",
  1895 => x"f5c282e8",
  1896 => x"807548ed",
  1897 => x"976e7e70",
  1898 => x"4b494bbf",
  1899 => x"a3c1486e",
  1900 => x"11816a50",
  1901 => x"58a6cc48",
  1902 => x"c402ac70",
  1903 => x"c0486e87",
  1904 => x"0566c850",
  1905 => x"f5c287c7",
  1906 => x"a5c448f1",
  1907 => x"c485c178",
  1908 => x"ff04adb7",
  1909 => x"dcc487c0",
  1910 => x"fdf5c287",
  1911 => x"b7c848bf",
  1912 => x"87d101a8",
  1913 => x"cc02acca",
  1914 => x"02accd87",
  1915 => x"b7c087c7",
  1916 => x"f3c003ac",
  1917 => x"fdf5c287",
  1918 => x"b7c84bbf",
  1919 => x"87d203ab",
  1920 => x"49c1f6c2",
  1921 => x"e0c08173",
  1922 => x"c883c151",
  1923 => x"ff04abb7",
  1924 => x"f6c287ee",
  1925 => x"d2c148c9",
  1926 => x"50cfc150",
  1927 => x"c050cdc1",
  1928 => x"c380e450",
  1929 => x"87cdc378",
  1930 => x"bffdf5c2",
  1931 => x"80c14849",
  1932 => x"58c1f6c2",
  1933 => x"81a0c448",
  1934 => x"f8c25174",
  1935 => x"b7f0c087",
  1936 => x"87da04ac",
  1937 => x"acb7f9c0",
  1938 => x"c287d301",
  1939 => x"49bff5f5",
  1940 => x"4a7491ca",
  1941 => x"c28af0c0",
  1942 => x"7248f5f5",
  1943 => x"acca78a1",
  1944 => x"87c6c002",
  1945 => x"c205accd",
  1946 => x"f5c287cb",
  1947 => x"78c348f1",
  1948 => x"c087c2c2",
  1949 => x"04acb7f0",
  1950 => x"f9c087db",
  1951 => x"c001acb7",
  1952 => x"f5c287d3",
  1953 => x"d049bff9",
  1954 => x"c04a7491",
  1955 => x"f5c28af0",
  1956 => x"a17248f9",
  1957 => x"b7c1c178",
  1958 => x"dbc004ac",
  1959 => x"b7c6c187",
  1960 => x"d3c001ac",
  1961 => x"f9f5c287",
  1962 => x"91d049bf",
  1963 => x"f7c04a74",
  1964 => x"f9f5c28a",
  1965 => x"78a17248",
  1966 => x"c002acca",
  1967 => x"accd87c6",
  1968 => x"87f1c005",
  1969 => x"48f1f5c2",
  1970 => x"e8c078c3",
  1971 => x"ace2c087",
  1972 => x"87c9c005",
  1973 => x"c048a6c4",
  1974 => x"d8c078fb",
  1975 => x"02acca87",
  1976 => x"cd87c6c0",
  1977 => x"c9c005ac",
  1978 => x"f1f5c287",
  1979 => x"c078c348",
  1980 => x"a6c887c3",
  1981 => x"acb7c05c",
  1982 => x"87c4c003",
  1983 => x"87cac048",
  1984 => x"f90266c4",
  1985 => x"c34887c6",
  1986 => x"8ef499ff",
  1987 => x"4387cff8",
  1988 => x"3d464e4f",
  1989 => x"444f4d00",
  1990 => x"4d414e00",
  1991 => x"45440045",
  1992 => x"4c554146",
  1993 => x"00303d54",
  1994 => x"00001f0f",
  1995 => x"00001f15",
  1996 => x"00001f19",
  1997 => x"00001f1e",
  1998 => x"48d0ff1e",
  1999 => x"7178c9c8",
  2000 => x"08d4ff48",
  2001 => x"1e4f2678",
  2002 => x"eb494a71",
  2003 => x"48d0ff87",
  2004 => x"4f2678c8",
  2005 => x"711e731e",
  2006 => x"d9f6c24b",
  2007 => x"87c302bf",
  2008 => x"ff87ebc2",
  2009 => x"c9c848d0",
  2010 => x"c0497378",
  2011 => x"d4ffb1e0",
  2012 => x"c2787148",
  2013 => x"c048cdf6",
  2014 => x"0266c878",
  2015 => x"ffc387c5",
  2016 => x"c087c249",
  2017 => x"d5f6c249",
  2018 => x"0266cc59",
  2019 => x"d5c587c6",
  2020 => x"87c44ad5",
  2021 => x"4affffcf",
  2022 => x"5ad9f6c2",
  2023 => x"48d9f6c2",
  2024 => x"87c478c1",
  2025 => x"4c264d26",
  2026 => x"4f264b26",
  2027 => x"5c5b5e0e",
  2028 => x"4a710e5d",
  2029 => x"bfd5f6c2",
  2030 => x"029a724c",
  2031 => x"c84987cb",
  2032 => x"cafdc191",
  2033 => x"c483714b",
  2034 => x"cac1c287",
  2035 => x"134dc04b",
  2036 => x"c2997449",
  2037 => x"b9bfd1f6",
  2038 => x"7148d4ff",
  2039 => x"2cb7c178",
  2040 => x"adb7c885",
  2041 => x"c287e804",
  2042 => x"48bfcdf6",
  2043 => x"f6c280c8",
  2044 => x"effe58d1",
  2045 => x"1e731e87",
  2046 => x"4a134b71",
  2047 => x"87cb029a",
  2048 => x"e7fe4972",
  2049 => x"9a4a1387",
  2050 => x"fe87f505",
  2051 => x"c21e87da",
  2052 => x"49bfcdf6",
  2053 => x"48cdf6c2",
  2054 => x"c478a1c1",
  2055 => x"03a9b7c0",
  2056 => x"d4ff87db",
  2057 => x"d1f6c248",
  2058 => x"f6c278bf",
  2059 => x"c249bfcd",
  2060 => x"c148cdf6",
  2061 => x"c0c478a1",
  2062 => x"e504a9b7",
  2063 => x"48d0ff87",
  2064 => x"f6c278c8",
  2065 => x"78c048d9",
  2066 => x"00004f26",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"005f5f00",
  2070 => x"03000000",
  2071 => x"03030003",
  2072 => x"7f140000",
  2073 => x"7f7f147f",
  2074 => x"24000014",
  2075 => x"3a6b6b2e",
  2076 => x"6a4c0012",
  2077 => x"566c1836",
  2078 => x"7e300032",
  2079 => x"3a77594f",
  2080 => x"00004068",
  2081 => x"00030704",
  2082 => x"00000000",
  2083 => x"41633e1c",
  2084 => x"00000000",
  2085 => x"1c3e6341",
  2086 => x"2a080000",
  2087 => x"3e1c1c3e",
  2088 => x"0800082a",
  2089 => x"083e3e08",
  2090 => x"00000008",
  2091 => x"0060e080",
  2092 => x"08000000",
  2093 => x"08080808",
  2094 => x"00000008",
  2095 => x"00606000",
  2096 => x"60400000",
  2097 => x"060c1830",
  2098 => x"3e000103",
  2099 => x"7f4d597f",
  2100 => x"0400003e",
  2101 => x"007f7f06",
  2102 => x"42000000",
  2103 => x"4f597163",
  2104 => x"22000046",
  2105 => x"7f494963",
  2106 => x"1c180036",
  2107 => x"7f7f1316",
  2108 => x"27000010",
  2109 => x"7d454567",
  2110 => x"3c000039",
  2111 => x"79494b7e",
  2112 => x"01000030",
  2113 => x"0f797101",
  2114 => x"36000007",
  2115 => x"7f49497f",
  2116 => x"06000036",
  2117 => x"3f69494f",
  2118 => x"0000001e",
  2119 => x"00666600",
  2120 => x"00000000",
  2121 => x"0066e680",
  2122 => x"08000000",
  2123 => x"22141408",
  2124 => x"14000022",
  2125 => x"14141414",
  2126 => x"22000014",
  2127 => x"08141422",
  2128 => x"02000008",
  2129 => x"0f595103",
  2130 => x"7f3e0006",
  2131 => x"1f555d41",
  2132 => x"7e00001e",
  2133 => x"7f09097f",
  2134 => x"7f00007e",
  2135 => x"7f49497f",
  2136 => x"1c000036",
  2137 => x"4141633e",
  2138 => x"7f000041",
  2139 => x"3e63417f",
  2140 => x"7f00001c",
  2141 => x"4149497f",
  2142 => x"7f000041",
  2143 => x"0109097f",
  2144 => x"3e000001",
  2145 => x"7b49417f",
  2146 => x"7f00007a",
  2147 => x"7f08087f",
  2148 => x"0000007f",
  2149 => x"417f7f41",
  2150 => x"20000000",
  2151 => x"7f404060",
  2152 => x"7f7f003f",
  2153 => x"63361c08",
  2154 => x"7f000041",
  2155 => x"4040407f",
  2156 => x"7f7f0040",
  2157 => x"7f060c06",
  2158 => x"7f7f007f",
  2159 => x"7f180c06",
  2160 => x"3e00007f",
  2161 => x"7f41417f",
  2162 => x"7f00003e",
  2163 => x"0f09097f",
  2164 => x"7f3e0006",
  2165 => x"7e7f6141",
  2166 => x"7f000040",
  2167 => x"7f19097f",
  2168 => x"26000066",
  2169 => x"7b594d6f",
  2170 => x"01000032",
  2171 => x"017f7f01",
  2172 => x"3f000001",
  2173 => x"7f40407f",
  2174 => x"0f00003f",
  2175 => x"3f70703f",
  2176 => x"7f7f000f",
  2177 => x"7f301830",
  2178 => x"6341007f",
  2179 => x"361c1c36",
  2180 => x"03014163",
  2181 => x"067c7c06",
  2182 => x"71610103",
  2183 => x"43474d59",
  2184 => x"00000041",
  2185 => x"41417f7f",
  2186 => x"03010000",
  2187 => x"30180c06",
  2188 => x"00004060",
  2189 => x"7f7f4141",
  2190 => x"0c080000",
  2191 => x"0c060306",
  2192 => x"80800008",
  2193 => x"80808080",
  2194 => x"00000080",
  2195 => x"04070300",
  2196 => x"20000000",
  2197 => x"7c545474",
  2198 => x"7f000078",
  2199 => x"7c44447f",
  2200 => x"38000038",
  2201 => x"4444447c",
  2202 => x"38000000",
  2203 => x"7f44447c",
  2204 => x"3800007f",
  2205 => x"5c54547c",
  2206 => x"04000018",
  2207 => x"05057f7e",
  2208 => x"18000000",
  2209 => x"fca4a4bc",
  2210 => x"7f00007c",
  2211 => x"7c04047f",
  2212 => x"00000078",
  2213 => x"407d3d00",
  2214 => x"80000000",
  2215 => x"7dfd8080",
  2216 => x"7f000000",
  2217 => x"6c38107f",
  2218 => x"00000044",
  2219 => x"407f3f00",
  2220 => x"7c7c0000",
  2221 => x"7c0c180c",
  2222 => x"7c000078",
  2223 => x"7c04047c",
  2224 => x"38000078",
  2225 => x"7c44447c",
  2226 => x"fc000038",
  2227 => x"3c2424fc",
  2228 => x"18000018",
  2229 => x"fc24243c",
  2230 => x"7c0000fc",
  2231 => x"0c04047c",
  2232 => x"48000008",
  2233 => x"7454545c",
  2234 => x"04000020",
  2235 => x"44447f3f",
  2236 => x"3c000000",
  2237 => x"7c40407c",
  2238 => x"1c00007c",
  2239 => x"3c60603c",
  2240 => x"7c3c001c",
  2241 => x"7c603060",
  2242 => x"6c44003c",
  2243 => x"6c381038",
  2244 => x"1c000044",
  2245 => x"3c60e0bc",
  2246 => x"4400001c",
  2247 => x"4c5c7464",
  2248 => x"08000044",
  2249 => x"41773e08",
  2250 => x"00000041",
  2251 => x"007f7f00",
  2252 => x"41000000",
  2253 => x"083e7741",
  2254 => x"01020008",
  2255 => x"02020301",
  2256 => x"7f7f0001",
  2257 => x"7f7f7f7f",
  2258 => x"0808007f",
  2259 => x"3e3e1c1c",
  2260 => x"7f7f7f7f",
  2261 => x"1c1c3e3e",
  2262 => x"10000808",
  2263 => x"187c7c18",
  2264 => x"10000010",
  2265 => x"307c7c30",
  2266 => x"30100010",
  2267 => x"1e786060",
  2268 => x"66420006",
  2269 => x"663c183c",
  2270 => x"38780042",
  2271 => x"6cc6c26a",
  2272 => x"00600038",
  2273 => x"00006000",
  2274 => x"5e0e0060",
  2275 => x"0e5d5c5b",
  2276 => x"c24c711e",
  2277 => x"4dbfeaf6",
  2278 => x"1ec04bc0",
  2279 => x"c702ab74",
  2280 => x"48a6c487",
  2281 => x"87c578c0",
  2282 => x"c148a6c4",
  2283 => x"1e66c478",
  2284 => x"dfee4973",
  2285 => x"c086c887",
  2286 => x"efef49e0",
  2287 => x"4aa5c487",
  2288 => x"f0f0496a",
  2289 => x"87c6f187",
  2290 => x"83c185cb",
  2291 => x"04abb7c8",
  2292 => x"2687c7ff",
  2293 => x"4c264d26",
  2294 => x"4f264b26",
  2295 => x"c24a711e",
  2296 => x"c25aeef6",
  2297 => x"c748eef6",
  2298 => x"ddfe4978",
  2299 => x"1e4f2687",
  2300 => x"4a711e73",
  2301 => x"03aab7c0",
  2302 => x"ddc287d3",
  2303 => x"c405bfcf",
  2304 => x"c24bc187",
  2305 => x"c24bc087",
  2306 => x"c45bd3dd",
  2307 => x"d3ddc287",
  2308 => x"cfddc25a",
  2309 => x"9ac14abf",
  2310 => x"49a2c0c1",
  2311 => x"fc87e8ec",
  2312 => x"cfddc248",
  2313 => x"effe78bf",
  2314 => x"4a711e87",
  2315 => x"721e66c4",
  2316 => x"dadfff49",
  2317 => x"4f262687",
  2318 => x"cfddc21e",
  2319 => x"dcff49bf",
  2320 => x"f6c287c2",
  2321 => x"bfe848e2",
  2322 => x"def6c278",
  2323 => x"78bfec48",
  2324 => x"bfe2f6c2",
  2325 => x"ffc3494a",
  2326 => x"2ab7c899",
  2327 => x"b0714872",
  2328 => x"58eaf6c2",
  2329 => x"5e0e4f26",
  2330 => x"0e5d5c5b",
  2331 => x"c7ff4b71",
  2332 => x"ddf6c287",
  2333 => x"7350c048",
  2334 => x"e7dbff49",
  2335 => x"4c497087",
  2336 => x"eecb9cc2",
  2337 => x"87cfcb49",
  2338 => x"c24d4970",
  2339 => x"bf97ddf6",
  2340 => x"87e4c105",
  2341 => x"c24966d0",
  2342 => x"99bfe6f6",
  2343 => x"d487d705",
  2344 => x"f6c24966",
  2345 => x"0599bfde",
  2346 => x"497387cc",
  2347 => x"87f4daff",
  2348 => x"c1029870",
  2349 => x"4cc187c2",
  2350 => x"7587fdfd",
  2351 => x"87e3ca49",
  2352 => x"c6029870",
  2353 => x"ddf6c287",
  2354 => x"c250c148",
  2355 => x"bf97ddf6",
  2356 => x"87e4c005",
  2357 => x"bfe6f6c2",
  2358 => x"9966d049",
  2359 => x"87d6ff05",
  2360 => x"bfdef6c2",
  2361 => x"9966d449",
  2362 => x"87caff05",
  2363 => x"d9ff4973",
  2364 => x"987087f2",
  2365 => x"87fefe05",
  2366 => x"d7fb4874",
  2367 => x"5b5e0e87",
  2368 => x"f40e5d5c",
  2369 => x"4c4dc086",
  2370 => x"c47ebfec",
  2371 => x"f6c248a6",
  2372 => x"c178bfea",
  2373 => x"c71ec01e",
  2374 => x"87cafd49",
  2375 => x"987086c8",
  2376 => x"ff87ce02",
  2377 => x"87c7fb49",
  2378 => x"ff49dac1",
  2379 => x"c187f5d8",
  2380 => x"ddf6c24d",
  2381 => x"c302bf97",
  2382 => x"87f9cd87",
  2383 => x"bfe2f6c2",
  2384 => x"cfddc24b",
  2385 => x"ebc005bf",
  2386 => x"49fdc387",
  2387 => x"87d4d8ff",
  2388 => x"ff49fac3",
  2389 => x"7387cdd8",
  2390 => x"99ffc349",
  2391 => x"49c01e71",
  2392 => x"7387c6fb",
  2393 => x"29b7c849",
  2394 => x"49c11e71",
  2395 => x"c887fafa",
  2396 => x"87c1c686",
  2397 => x"bfe6f6c2",
  2398 => x"dd029b4b",
  2399 => x"cbddc287",
  2400 => x"dec749bf",
  2401 => x"05987087",
  2402 => x"4bc087c4",
  2403 => x"e0c287d2",
  2404 => x"87c3c749",
  2405 => x"58cfddc2",
  2406 => x"ddc287c6",
  2407 => x"78c048cb",
  2408 => x"99c24973",
  2409 => x"c387ce05",
  2410 => x"d6ff49eb",
  2411 => x"497087f6",
  2412 => x"c20299c2",
  2413 => x"734cfb87",
  2414 => x"0599c149",
  2415 => x"f4c387ce",
  2416 => x"dfd6ff49",
  2417 => x"c2497087",
  2418 => x"87c20299",
  2419 => x"49734cfa",
  2420 => x"ce0599c8",
  2421 => x"49f5c387",
  2422 => x"87c8d6ff",
  2423 => x"99c24970",
  2424 => x"c287d502",
  2425 => x"02bfeef6",
  2426 => x"c14887ca",
  2427 => x"f2f6c288",
  2428 => x"87c2c058",
  2429 => x"4dc14cff",
  2430 => x"99c44973",
  2431 => x"c387ce05",
  2432 => x"d5ff49f2",
  2433 => x"497087de",
  2434 => x"dc0299c2",
  2435 => x"eef6c287",
  2436 => x"c7487ebf",
  2437 => x"c003a8b7",
  2438 => x"486e87cb",
  2439 => x"f6c280c1",
  2440 => x"c2c058f2",
  2441 => x"c14cfe87",
  2442 => x"49fdc34d",
  2443 => x"87f4d4ff",
  2444 => x"99c24970",
  2445 => x"87d5c002",
  2446 => x"bfeef6c2",
  2447 => x"87c9c002",
  2448 => x"48eef6c2",
  2449 => x"c2c078c0",
  2450 => x"c14cfd87",
  2451 => x"49fac34d",
  2452 => x"87d0d4ff",
  2453 => x"99c24970",
  2454 => x"87d9c002",
  2455 => x"bfeef6c2",
  2456 => x"a8b7c748",
  2457 => x"87c9c003",
  2458 => x"48eef6c2",
  2459 => x"c2c078c7",
  2460 => x"c14cfc87",
  2461 => x"acb7c04d",
  2462 => x"87d1c003",
  2463 => x"c14a66c4",
  2464 => x"026a82d8",
  2465 => x"6a87c6c0",
  2466 => x"7349744b",
  2467 => x"c31ec00f",
  2468 => x"dac11ef0",
  2469 => x"87cef749",
  2470 => x"987086c8",
  2471 => x"87e2c002",
  2472 => x"c248a6c8",
  2473 => x"78bfeef6",
  2474 => x"cb4966c8",
  2475 => x"4866c491",
  2476 => x"7e708071",
  2477 => x"c002bf6e",
  2478 => x"bf6e87c8",
  2479 => x"4966c84b",
  2480 => x"9d750f73",
  2481 => x"87c8c002",
  2482 => x"bfeef6c2",
  2483 => x"87faf249",
  2484 => x"bfd3ddc2",
  2485 => x"87ddc002",
  2486 => x"87c7c249",
  2487 => x"c0029870",
  2488 => x"f6c287d3",
  2489 => x"f249bfee",
  2490 => x"49c087e0",
  2491 => x"c287c0f4",
  2492 => x"c048d3dd",
  2493 => x"f38ef478",
  2494 => x"5e0e87da",
  2495 => x"0e5d5c5b",
  2496 => x"c24c711e",
  2497 => x"49bfeaf6",
  2498 => x"4da1cdc1",
  2499 => x"6981d1c1",
  2500 => x"029c747e",
  2501 => x"a5c487cf",
  2502 => x"c27b744b",
  2503 => x"49bfeaf6",
  2504 => x"6e87f9f2",
  2505 => x"059c747b",
  2506 => x"4bc087c4",
  2507 => x"4bc187c2",
  2508 => x"faf24973",
  2509 => x"0266d487",
  2510 => x"da4987c7",
  2511 => x"c24a7087",
  2512 => x"c24ac087",
  2513 => x"265ad7dd",
  2514 => x"0087c9f2",
  2515 => x"00000000",
  2516 => x"00000000",
  2517 => x"1e000000",
  2518 => x"c8ff4a71",
  2519 => x"a17249bf",
  2520 => x"1e4f2648",
  2521 => x"89bfc8ff",
  2522 => x"c0c0c0fe",
  2523 => x"01a9c0c0",
  2524 => x"4ac087c4",
  2525 => x"4ac187c2",
  2526 => x"4f264872",
  2527 => x"5c5b5e0e",
  2528 => x"711e0e5d",
  2529 => x"4bd4ff4d",
  2530 => x"f6c21e75",
  2531 => x"c1fe49f2",
  2532 => x"86c487d0",
  2533 => x"026e7e70",
  2534 => x"c287ffc3",
  2535 => x"4cbffaf6",
  2536 => x"dafe4975",
  2537 => x"a8de87fe",
  2538 => x"87ebc005",
  2539 => x"d3ff4975",
  2540 => x"987087ec",
  2541 => x"c287db02",
  2542 => x"1ebff5f5",
  2543 => x"ff49e1c0",
  2544 => x"c487f7d0",
  2545 => x"f4e2c286",
  2546 => x"c250c048",
  2547 => x"fe49c1f6",
  2548 => x"48c187ea",
  2549 => x"ff87c5c3",
  2550 => x"c5c848d0",
  2551 => x"7bd6c178",
  2552 => x"976e4ac0",
  2553 => x"486e7bbf",
  2554 => x"7e7080c1",
  2555 => x"e0c082c1",
  2556 => x"ff04aab7",
  2557 => x"d0ff87ec",
  2558 => x"c878c448",
  2559 => x"d3c178c5",
  2560 => x"c47bc17b",
  2561 => x"029c7478",
  2562 => x"c287fdc1",
  2563 => x"c87eeee4",
  2564 => x"c08c4dc0",
  2565 => x"c603acb7",
  2566 => x"a4c0c887",
  2567 => x"c24cc04d",
  2568 => x"bf97dff1",
  2569 => x"0299d049",
  2570 => x"1ec087d2",
  2571 => x"49f2f6c2",
  2572 => x"87cac2fe",
  2573 => x"497086c4",
  2574 => x"87efc04a",
  2575 => x"1eeee4c2",
  2576 => x"49f2f6c2",
  2577 => x"87f6c1fe",
  2578 => x"497086c4",
  2579 => x"48d0ff4a",
  2580 => x"c178c5c8",
  2581 => x"976e7bd4",
  2582 => x"486e7bbf",
  2583 => x"7e7080c1",
  2584 => x"ff058dc1",
  2585 => x"d0ff87f0",
  2586 => x"7278c448",
  2587 => x"c5c0059a",
  2588 => x"c048c087",
  2589 => x"1ec187e6",
  2590 => x"49f2f6c2",
  2591 => x"87ddfffd",
  2592 => x"9c7486c4",
  2593 => x"87c3fe05",
  2594 => x"c848d0ff",
  2595 => x"d3c178c5",
  2596 => x"c47bc07b",
  2597 => x"c048c178",
  2598 => x"48c087c2",
  2599 => x"264d2626",
  2600 => x"264b264c",
  2601 => x"4a711e4f",
  2602 => x"c50566c4",
  2603 => x"fb497287",
  2604 => x"4f2687ca",
  2605 => x"e4c21e00",
  2606 => x"c149bfc3",
  2607 => x"c7e4c2b9",
  2608 => x"48d4ff59",
  2609 => x"ff78ffc3",
  2610 => x"e1c848d0",
  2611 => x"48d4ff78",
  2612 => x"31c478c1",
  2613 => x"d0ff7871",
  2614 => x"78e0c048",
  2615 => x"c21e4f26",
  2616 => x"c21ef7e3",
  2617 => x"fd49f2f6",
  2618 => x"c487f7fb",
  2619 => x"02987086",
  2620 => x"c0ff87c3",
  2621 => x"314f2687",
  2622 => x"5a484b35",
  2623 => x"43202020",
  2624 => x"00004746",
  2625 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
