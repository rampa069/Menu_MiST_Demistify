library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"e7fe4972",
     1 => x"9a4a1387",
     2 => x"fe87f505",
     3 => x"c21e87da",
     4 => x"49bfcdf6",
     5 => x"48cdf6c2",
     6 => x"c478a1c1",
     7 => x"03a9b7c0",
     8 => x"d4ff87db",
     9 => x"d1f6c248",
    10 => x"f6c278bf",
    11 => x"c249bfcd",
    12 => x"c148cdf6",
    13 => x"c0c478a1",
    14 => x"e504a9b7",
    15 => x"48d0ff87",
    16 => x"f6c278c8",
    17 => x"78c048d9",
    18 => x"00004f26",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"005f5f00",
    22 => x"03000000",
    23 => x"03030003",
    24 => x"7f140000",
    25 => x"7f7f147f",
    26 => x"24000014",
    27 => x"3a6b6b2e",
    28 => x"6a4c0012",
    29 => x"566c1836",
    30 => x"7e300032",
    31 => x"3a77594f",
    32 => x"00004068",
    33 => x"00030704",
    34 => x"00000000",
    35 => x"41633e1c",
    36 => x"00000000",
    37 => x"1c3e6341",
    38 => x"2a080000",
    39 => x"3e1c1c3e",
    40 => x"0800082a",
    41 => x"083e3e08",
    42 => x"00000008",
    43 => x"0060e080",
    44 => x"08000000",
    45 => x"08080808",
    46 => x"00000008",
    47 => x"00606000",
    48 => x"60400000",
    49 => x"060c1830",
    50 => x"3e000103",
    51 => x"7f4d597f",
    52 => x"0400003e",
    53 => x"007f7f06",
    54 => x"42000000",
    55 => x"4f597163",
    56 => x"22000046",
    57 => x"7f494963",
    58 => x"1c180036",
    59 => x"7f7f1316",
    60 => x"27000010",
    61 => x"7d454567",
    62 => x"3c000039",
    63 => x"79494b7e",
    64 => x"01000030",
    65 => x"0f797101",
    66 => x"36000007",
    67 => x"7f49497f",
    68 => x"06000036",
    69 => x"3f69494f",
    70 => x"0000001e",
    71 => x"00666600",
    72 => x"00000000",
    73 => x"0066e680",
    74 => x"08000000",
    75 => x"22141408",
    76 => x"14000022",
    77 => x"14141414",
    78 => x"22000014",
    79 => x"08141422",
    80 => x"02000008",
    81 => x"0f595103",
    82 => x"7f3e0006",
    83 => x"1f555d41",
    84 => x"7e00001e",
    85 => x"7f09097f",
    86 => x"7f00007e",
    87 => x"7f49497f",
    88 => x"1c000036",
    89 => x"4141633e",
    90 => x"7f000041",
    91 => x"3e63417f",
    92 => x"7f00001c",
    93 => x"4149497f",
    94 => x"7f000041",
    95 => x"0109097f",
    96 => x"3e000001",
    97 => x"7b49417f",
    98 => x"7f00007a",
    99 => x"7f08087f",
   100 => x"0000007f",
   101 => x"417f7f41",
   102 => x"20000000",
   103 => x"7f404060",
   104 => x"7f7f003f",
   105 => x"63361c08",
   106 => x"7f000041",
   107 => x"4040407f",
   108 => x"7f7f0040",
   109 => x"7f060c06",
   110 => x"7f7f007f",
   111 => x"7f180c06",
   112 => x"3e00007f",
   113 => x"7f41417f",
   114 => x"7f00003e",
   115 => x"0f09097f",
   116 => x"7f3e0006",
   117 => x"7e7f6141",
   118 => x"7f000040",
   119 => x"7f19097f",
   120 => x"26000066",
   121 => x"7b594d6f",
   122 => x"01000032",
   123 => x"017f7f01",
   124 => x"3f000001",
   125 => x"7f40407f",
   126 => x"0f00003f",
   127 => x"3f70703f",
   128 => x"7f7f000f",
   129 => x"7f301830",
   130 => x"6341007f",
   131 => x"361c1c36",
   132 => x"03014163",
   133 => x"067c7c06",
   134 => x"71610103",
   135 => x"43474d59",
   136 => x"00000041",
   137 => x"41417f7f",
   138 => x"03010000",
   139 => x"30180c06",
   140 => x"00004060",
   141 => x"7f7f4141",
   142 => x"0c080000",
   143 => x"0c060306",
   144 => x"80800008",
   145 => x"80808080",
   146 => x"00000080",
   147 => x"04070300",
   148 => x"20000000",
   149 => x"7c545474",
   150 => x"7f000078",
   151 => x"7c44447f",
   152 => x"38000038",
   153 => x"4444447c",
   154 => x"38000000",
   155 => x"7f44447c",
   156 => x"3800007f",
   157 => x"5c54547c",
   158 => x"04000018",
   159 => x"05057f7e",
   160 => x"18000000",
   161 => x"fca4a4bc",
   162 => x"7f00007c",
   163 => x"7c04047f",
   164 => x"00000078",
   165 => x"407d3d00",
   166 => x"80000000",
   167 => x"7dfd8080",
   168 => x"7f000000",
   169 => x"6c38107f",
   170 => x"00000044",
   171 => x"407f3f00",
   172 => x"7c7c0000",
   173 => x"7c0c180c",
   174 => x"7c000078",
   175 => x"7c04047c",
   176 => x"38000078",
   177 => x"7c44447c",
   178 => x"fc000038",
   179 => x"3c2424fc",
   180 => x"18000018",
   181 => x"fc24243c",
   182 => x"7c0000fc",
   183 => x"0c04047c",
   184 => x"48000008",
   185 => x"7454545c",
   186 => x"04000020",
   187 => x"44447f3f",
   188 => x"3c000000",
   189 => x"7c40407c",
   190 => x"1c00007c",
   191 => x"3c60603c",
   192 => x"7c3c001c",
   193 => x"7c603060",
   194 => x"6c44003c",
   195 => x"6c381038",
   196 => x"1c000044",
   197 => x"3c60e0bc",
   198 => x"4400001c",
   199 => x"4c5c7464",
   200 => x"08000044",
   201 => x"41773e08",
   202 => x"00000041",
   203 => x"007f7f00",
   204 => x"41000000",
   205 => x"083e7741",
   206 => x"01020008",
   207 => x"02020301",
   208 => x"7f7f0001",
   209 => x"7f7f7f7f",
   210 => x"0808007f",
   211 => x"3e3e1c1c",
   212 => x"7f7f7f7f",
   213 => x"1c1c3e3e",
   214 => x"10000808",
   215 => x"187c7c18",
   216 => x"10000010",
   217 => x"307c7c30",
   218 => x"30100010",
   219 => x"1e786060",
   220 => x"66420006",
   221 => x"663c183c",
   222 => x"38780042",
   223 => x"6cc6c26a",
   224 => x"00600038",
   225 => x"00006000",
   226 => x"5e0e0060",
   227 => x"0e5d5c5b",
   228 => x"c24c711e",
   229 => x"4dbfeaf6",
   230 => x"1ec04bc0",
   231 => x"c702ab74",
   232 => x"48a6c487",
   233 => x"87c578c0",
   234 => x"c148a6c4",
   235 => x"1e66c478",
   236 => x"dfee4973",
   237 => x"c086c887",
   238 => x"efef49e0",
   239 => x"4aa5c487",
   240 => x"f0f0496a",
   241 => x"87c6f187",
   242 => x"83c185cb",
   243 => x"04abb7c8",
   244 => x"2687c7ff",
   245 => x"4c264d26",
   246 => x"4f264b26",
   247 => x"c24a711e",
   248 => x"c25aeef6",
   249 => x"c748eef6",
   250 => x"ddfe4978",
   251 => x"1e4f2687",
   252 => x"4a711e73",
   253 => x"03aab7c0",
   254 => x"ddc287d3",
   255 => x"c405bfcf",
   256 => x"c24bc187",
   257 => x"c24bc087",
   258 => x"c45bd3dd",
   259 => x"d3ddc287",
   260 => x"cfddc25a",
   261 => x"9ac14abf",
   262 => x"49a2c0c1",
   263 => x"fc87e8ec",
   264 => x"cfddc248",
   265 => x"effe78bf",
   266 => x"4a711e87",
   267 => x"721e66c4",
   268 => x"dadfff49",
   269 => x"4f262687",
   270 => x"cfddc21e",
   271 => x"dcff49bf",
   272 => x"f6c287c2",
   273 => x"bfe848e2",
   274 => x"def6c278",
   275 => x"78bfec48",
   276 => x"bfe2f6c2",
   277 => x"ffc3494a",
   278 => x"2ab7c899",
   279 => x"b0714872",
   280 => x"58eaf6c2",
   281 => x"5e0e4f26",
   282 => x"0e5d5c5b",
   283 => x"c7ff4b71",
   284 => x"ddf6c287",
   285 => x"7350c048",
   286 => x"e7dbff49",
   287 => x"4c497087",
   288 => x"eecb9cc2",
   289 => x"87cfcb49",
   290 => x"c24d4970",
   291 => x"bf97ddf6",
   292 => x"87e4c105",
   293 => x"c24966d0",
   294 => x"99bfe6f6",
   295 => x"d487d705",
   296 => x"f6c24966",
   297 => x"0599bfde",
   298 => x"497387cc",
   299 => x"87f4daff",
   300 => x"c1029870",
   301 => x"4cc187c2",
   302 => x"7587fdfd",
   303 => x"87e3ca49",
   304 => x"c6029870",
   305 => x"ddf6c287",
   306 => x"c250c148",
   307 => x"bf97ddf6",
   308 => x"87e4c005",
   309 => x"bfe6f6c2",
   310 => x"9966d049",
   311 => x"87d6ff05",
   312 => x"bfdef6c2",
   313 => x"9966d449",
   314 => x"87caff05",
   315 => x"d9ff4973",
   316 => x"987087f2",
   317 => x"87fefe05",
   318 => x"d7fb4874",
   319 => x"5b5e0e87",
   320 => x"f40e5d5c",
   321 => x"4c4dc086",
   322 => x"c47ebfec",
   323 => x"f6c248a6",
   324 => x"c178bfea",
   325 => x"c71ec01e",
   326 => x"87cafd49",
   327 => x"987086c8",
   328 => x"ff87ce02",
   329 => x"87c7fb49",
   330 => x"ff49dac1",
   331 => x"c187f5d8",
   332 => x"ddf6c24d",
   333 => x"c302bf97",
   334 => x"87f9cd87",
   335 => x"bfe2f6c2",
   336 => x"cfddc24b",
   337 => x"ebc005bf",
   338 => x"49fdc387",
   339 => x"87d4d8ff",
   340 => x"ff49fac3",
   341 => x"7387cdd8",
   342 => x"99ffc349",
   343 => x"49c01e71",
   344 => x"7387c6fb",
   345 => x"29b7c849",
   346 => x"49c11e71",
   347 => x"c887fafa",
   348 => x"87c1c686",
   349 => x"bfe6f6c2",
   350 => x"dd029b4b",
   351 => x"cbddc287",
   352 => x"dec749bf",
   353 => x"05987087",
   354 => x"4bc087c4",
   355 => x"e0c287d2",
   356 => x"87c3c749",
   357 => x"58cfddc2",
   358 => x"ddc287c6",
   359 => x"78c048cb",
   360 => x"99c24973",
   361 => x"c387ce05",
   362 => x"d6ff49eb",
   363 => x"497087f6",
   364 => x"c20299c2",
   365 => x"734cfb87",
   366 => x"0599c149",
   367 => x"f4c387ce",
   368 => x"dfd6ff49",
   369 => x"c2497087",
   370 => x"87c20299",
   371 => x"49734cfa",
   372 => x"ce0599c8",
   373 => x"49f5c387",
   374 => x"87c8d6ff",
   375 => x"99c24970",
   376 => x"c287d502",
   377 => x"02bfeef6",
   378 => x"c14887ca",
   379 => x"f2f6c288",
   380 => x"87c2c058",
   381 => x"4dc14cff",
   382 => x"99c44973",
   383 => x"c387ce05",
   384 => x"d5ff49f2",
   385 => x"497087de",
   386 => x"dc0299c2",
   387 => x"eef6c287",
   388 => x"c7487ebf",
   389 => x"c003a8b7",
   390 => x"486e87cb",
   391 => x"f6c280c1",
   392 => x"c2c058f2",
   393 => x"c14cfe87",
   394 => x"49fdc34d",
   395 => x"87f4d4ff",
   396 => x"99c24970",
   397 => x"87d5c002",
   398 => x"bfeef6c2",
   399 => x"87c9c002",
   400 => x"48eef6c2",
   401 => x"c2c078c0",
   402 => x"c14cfd87",
   403 => x"49fac34d",
   404 => x"87d0d4ff",
   405 => x"99c24970",
   406 => x"87d9c002",
   407 => x"bfeef6c2",
   408 => x"a8b7c748",
   409 => x"87c9c003",
   410 => x"48eef6c2",
   411 => x"c2c078c7",
   412 => x"c14cfc87",
   413 => x"acb7c04d",
   414 => x"87d1c003",
   415 => x"c14a66c4",
   416 => x"026a82d8",
   417 => x"6a87c6c0",
   418 => x"7349744b",
   419 => x"c31ec00f",
   420 => x"dac11ef0",
   421 => x"87cef749",
   422 => x"987086c8",
   423 => x"87e2c002",
   424 => x"c248a6c8",
   425 => x"78bfeef6",
   426 => x"cb4966c8",
   427 => x"4866c491",
   428 => x"7e708071",
   429 => x"c002bf6e",
   430 => x"bf6e87c8",
   431 => x"4966c84b",
   432 => x"9d750f73",
   433 => x"87c8c002",
   434 => x"bfeef6c2",
   435 => x"87faf249",
   436 => x"bfd3ddc2",
   437 => x"87ddc002",
   438 => x"87c7c249",
   439 => x"c0029870",
   440 => x"f6c287d3",
   441 => x"f249bfee",
   442 => x"49c087e0",
   443 => x"c287c0f4",
   444 => x"c048d3dd",
   445 => x"f38ef478",
   446 => x"5e0e87da",
   447 => x"0e5d5c5b",
   448 => x"c24c711e",
   449 => x"49bfeaf6",
   450 => x"4da1cdc1",
   451 => x"6981d1c1",
   452 => x"029c747e",
   453 => x"a5c487cf",
   454 => x"c27b744b",
   455 => x"49bfeaf6",
   456 => x"6e87f9f2",
   457 => x"059c747b",
   458 => x"4bc087c4",
   459 => x"4bc187c2",
   460 => x"faf24973",
   461 => x"0266d487",
   462 => x"da4987c7",
   463 => x"c24a7087",
   464 => x"c24ac087",
   465 => x"265ad7dd",
   466 => x"0087c9f2",
   467 => x"00000000",
   468 => x"00000000",
   469 => x"1e000000",
   470 => x"c8ff4a71",
   471 => x"a17249bf",
   472 => x"1e4f2648",
   473 => x"89bfc8ff",
   474 => x"c0c0c0fe",
   475 => x"01a9c0c0",
   476 => x"4ac087c4",
   477 => x"4ac187c2",
   478 => x"4f264872",
   479 => x"5c5b5e0e",
   480 => x"711e0e5d",
   481 => x"4bd4ff4d",
   482 => x"f6c21e75",
   483 => x"c1fe49f2",
   484 => x"86c487d0",
   485 => x"026e7e70",
   486 => x"c287ffc3",
   487 => x"4cbffaf6",
   488 => x"dafe4975",
   489 => x"a8de87fe",
   490 => x"87ebc005",
   491 => x"d3ff4975",
   492 => x"987087ec",
   493 => x"c287db02",
   494 => x"1ebff5f5",
   495 => x"ff49e1c0",
   496 => x"c487f7d0",
   497 => x"f4e2c286",
   498 => x"c250c048",
   499 => x"fe49c1f6",
   500 => x"48c187ea",
   501 => x"ff87c5c3",
   502 => x"c5c848d0",
   503 => x"7bd6c178",
   504 => x"976e4ac0",
   505 => x"486e7bbf",
   506 => x"7e7080c1",
   507 => x"e0c082c1",
   508 => x"ff04aab7",
   509 => x"d0ff87ec",
   510 => x"c878c448",
   511 => x"d3c178c5",
   512 => x"c47bc17b",
   513 => x"029c7478",
   514 => x"c287fdc1",
   515 => x"c87eeee4",
   516 => x"c08c4dc0",
   517 => x"c603acb7",
   518 => x"a4c0c887",
   519 => x"c24cc04d",
   520 => x"bf97dff1",
   521 => x"0299d049",
   522 => x"1ec087d2",
   523 => x"49f2f6c2",
   524 => x"87cac2fe",
   525 => x"497086c4",
   526 => x"87efc04a",
   527 => x"1eeee4c2",
   528 => x"49f2f6c2",
   529 => x"87f6c1fe",
   530 => x"497086c4",
   531 => x"48d0ff4a",
   532 => x"c178c5c8",
   533 => x"976e7bd4",
   534 => x"486e7bbf",
   535 => x"7e7080c1",
   536 => x"ff058dc1",
   537 => x"d0ff87f0",
   538 => x"7278c448",
   539 => x"c5c0059a",
   540 => x"c048c087",
   541 => x"1ec187e6",
   542 => x"49f2f6c2",
   543 => x"87ddfffd",
   544 => x"9c7486c4",
   545 => x"87c3fe05",
   546 => x"c848d0ff",
   547 => x"d3c178c5",
   548 => x"c47bc07b",
   549 => x"c048c178",
   550 => x"48c087c2",
   551 => x"264d2626",
   552 => x"264b264c",
   553 => x"4a711e4f",
   554 => x"c50566c4",
   555 => x"fb497287",
   556 => x"4f2687ca",
   557 => x"e4c21e00",
   558 => x"c149bfc3",
   559 => x"c7e4c2b9",
   560 => x"48d4ff59",
   561 => x"ff78ffc3",
   562 => x"e1c848d0",
   563 => x"48d4ff78",
   564 => x"31c478c1",
   565 => x"d0ff7871",
   566 => x"78e0c048",
   567 => x"c21e4f26",
   568 => x"c21ef7e3",
   569 => x"fd49f2f6",
   570 => x"c487f7fb",
   571 => x"02987086",
   572 => x"c0ff87c3",
   573 => x"314f2687",
   574 => x"5a484b35",
   575 => x"43202020",
   576 => x"00004746",
   577 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
